// Verilog File 
module des (pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,pi133,pi134,pi135,pi136,pi137,pi138,
pi139,pi140,pi141,pi142,pi143,pi144,pi145,pi146,pi147,pi148,
pi149,pi150,pi151,pi152,pi153,pi154,pi155,pi156,pi157,pi158,
pi159,pi160,pi161,pi162,pi163,pi164,pi165,pi166,pi167,pi168,
pi169,pi170,pi171,pi172,pi173,pi174,pi175,pi176,pi177,pi178,
pi179,pi180,pi181,pi182,pi183,pi184,pi185,pi186,pi187,pi188,
pi189,pi190,pi191,pi192,pi193,pi194,pi195,pi196,pi197,pi198,
pi199,pi200,pi201,pi202,pi203,pi204,pi205,pi206,pi207,pi208,
pi209,pi210,pi211,pi212,pi213,pi214,pi215,pi216,pi217,pi218,
pi219,pi220,pi221,pi222,pi223,pi224,pi225,pi226,pi227,pi228,
pi229,pi230,pi231,pi232,pi233,pi234,pi235,pi236,pi237,pi238,
pi239,pi240,pi241,pi242,pi243,pi244,pi245,pi246,pi247,pi248,
pi249,pi250,pi251,pi252,pi253,pi254,pi255,po000,po001,po002,
po003,po004,po005,po006,po007,po008,po009,po010,po011,po012,
po013,po014,po015,po016,po017,po018,po019,po020,po021,po022,
po023,po024,po025,po026,po027,po028,po029,po030,po031,po032,
po033,po034,po035,po036,po037,po038,po039,po040,po041,po042,
po043,po044,po045,po046,po047,po048,po049,po050,po051,po052,
po053,po054,po055,po056,po057,po058,po059,po060,po061,po062,
po063,po064,po065,po066,po067,po068,po069,po070,po071,po072,
po073,po074,po075,po076,po077,po078,po079,po080,po081,po082,
po083,po084,po085,po086,po087,po088,po089,po090,po091,po092,
po093,po094,po095,po096,po097,po098,po099,po100,po101,po102,
po103,po104,po105,po106,po107,po108,po109,po110,po111,po112,
po113,po114,po115,po116,po117,po118,po119,po120,po121,po122,
po123,po124,po125,po126,po127,po128,po129,po130,po131,po132,
po133,po134,po135,po136,po137,po138,po139,po140,po141,po142,
po143,po144,po145,po146,po147,po148,po149,po150,po151,po152,
po153,po154,po155,po156,po157,po158,po159,po160,po161,po162,
po163,po164,po165,po166,po167,po168,po169,po170,po171,po172,
po173,po174,po175,po176,po177,po178,po179,po180,po181,po182,
po183,po184,po185,po186,po187,po188,po189,po190,po191,po192,
po193,po194,po195,po196,po197,po198,po199,po200,po201,po202,
po203,po204,po205,po206,po207,po208,po209,po210,po211,po212,
po213,po214,po215,po216,po217,po218,po219,po220,po221,po222,
po223,po224,po225,po226,po227,po228,po229,po230,po231,po232,
po233,po234,po235,po236,po237,po238,po239,po240,po241,po242,
po243,po244);

input pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,pi133,pi134,pi135,pi136,pi137,pi138,
pi139,pi140,pi141,pi142,pi143,pi144,pi145,pi146,pi147,pi148,
pi149,pi150,pi151,pi152,pi153,pi154,pi155,pi156,pi157,pi158,
pi159,pi160,pi161,pi162,pi163,pi164,pi165,pi166,pi167,pi168,
pi169,pi170,pi171,pi172,pi173,pi174,pi175,pi176,pi177,pi178,
pi179,pi180,pi181,pi182,pi183,pi184,pi185,pi186,pi187,pi188,
pi189,pi190,pi191,pi192,pi193,pi194,pi195,pi196,pi197,pi198,
pi199,pi200,pi201,pi202,pi203,pi204,pi205,pi206,pi207,pi208,
pi209,pi210,pi211,pi212,pi213,pi214,pi215,pi216,pi217,pi218,
pi219,pi220,pi221,pi222,pi223,pi224,pi225,pi226,pi227,pi228,
pi229,pi230,pi231,pi232,pi233,pi234,pi235,pi236,pi237,pi238,
pi239,pi240,pi241,pi242,pi243,pi244,pi245,pi246,pi247,pi248,
pi249,pi250,pi251,pi252,pi253,pi254,pi255;

output po000,po001,po002,po003,po004,po005,po006,po007,po008,
po009,po010,po011,po012,po013,po014,po015,po016,po017,po018,
po019,po020,po021,po022,po023,po024,po025,po026,po027,po028,
po029,po030,po031,po032,po033,po034,po035,po036,po037,po038,
po039,po040,po041,po042,po043,po044,po045,po046,po047,po048,
po049,po050,po051,po052,po053,po054,po055,po056,po057,po058,
po059,po060,po061,po062,po063,po064,po065,po066,po067,po068,
po069,po070,po071,po072,po073,po074,po075,po076,po077,po078,
po079,po080,po081,po082,po083,po084,po085,po086,po087,po088,
po089,po090,po091,po092,po093,po094,po095,po096,po097,po098,
po099,po100,po101,po102,po103,po104,po105,po106,po107,po108,
po109,po110,po111,po112,po113,po114,po115,po116,po117,po118,
po119,po120,po121,po122,po123,po124,po125,po126,po127,po128,
po129,po130,po131,po132,po133,po134,po135,po136,po137,po138,
po139,po140,po141,po142,po143,po144,po145,po146,po147,po148,
po149,po150,po151,po152,po153,po154,po155,po156,po157,po158,
po159,po160,po161,po162,po163,po164,po165,po166,po167,po168,
po169,po170,po171,po172,po173,po174,po175,po176,po177,po178,
po179,po180,po181,po182,po183,po184,po185,po186,po187,po188,
po189,po190,po191,po192,po193,po194,po195,po196,po197,po198,
po199,po200,po201,po202,po203,po204,po205,po206,po207,po208,
po209,po210,po211,po212,po213,po214,po215,po216,po217,po218,
po219,po220,po221,po222,po223,po224,po225,po226,po227,po228,
po229,po230,po231,po232,po233,po234,po235,po236,po237,po238,
po239,po240,po241,po242,po243,po244;

wire n501,n502,n503,n504,n505,n506,n507,n508,n509,
n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,
n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,
n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,
n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,
n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,
n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,
n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,
n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,
n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,
n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,
n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,
n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,
n630,n632,n633,n634,n635,n636,n637,n639,n640,n641,
n642,n643,n644,n646,n647,n648,n649,n650,n651,n653,
n654,n655,n656,n657,n658,n660,n661,n662,n663,n664,
n665,n667,n668,n669,n670,n671,n672,n674,n675,n676,
n677,n678,n679,n681,n682,n683,n684,n685,n686,n688,
n689,n690,n691,n692,n693,n695,n696,n697,n698,n699,
n700,n702,n703,n704,n705,n706,n707,n709,n710,n711,
n712,n713,n714,n716,n717,n718,n719,n720,n721,n723,
n724,n725,n726,n727,n728,n730,n731,n732,n733,n734,
n735,n737,n738,n739,n740,n741,n742,n744,n745,n746,
n747,n748,n749,n751,n752,n753,n754,n755,n756,n758,
n759,n760,n761,n762,n763,n765,n766,n767,n768,n769,
n770,n772,n773,n774,n775,n776,n777,n779,n780,n781,
n782,n783,n784,n786,n787,n788,n789,n790,n791,n793,
n794,n795,n796,n797,n798,n800,n801,n802,n803,n804,
n805,n807,n808,n809,n810,n811,n812,n814,n815,n816,
n817,n818,n819,n821,n822,n823,n824,n825,n826,n828,
n829,n830,n831,n832,n833,n835,n836,n837,n838,n839,
n840,n842,n843,n844,n845,n846,n847,n849,n850,n851,
n852,n853,n854,n856,n857,n858,n859,n860,n861,n863,
n864,n865,n866,n867,n868,n870,n871,n872,n873,n874,
n875,n877,n878,n879,n880,n881,n882,n884,n885,n886,
n887,n888,n889,n891,n892,n893,n894,n895,n896,n898,
n899,n900,n901,n902,n903,n905,n906,n907,n908,n909,
n910,n912,n913,n914,n915,n916,n917,n919,n920,n921,
n922,n923,n924,n926,n927,n928,n929,n930,n931,n933,
n934,n935,n936,n937,n938,n940,n941,n942,n943,n944,
n945,n947,n948,n949,n950,n951,n952,n954,n955,n956,
n957,n958,n959,n961,n962,n963,n964,n965,n966,n968,
n969,n970,n971,n972,n973,n975,n976,n977,n978,n979,
n980,n982,n983,n984,n985,n986,n987,n989,n990,n991,
n992,n993,n994,n996,n997,n998,n999,n1000,n1001,n1003,
n1004,n1005,n1006,n1007,n1008,n1010,n1011,n1012,n1013,n1014,
n1015,n1017,n1018,n1019,n1020,n1021,n1022,n1023,n1024,n1025,
n1026,n1027,n1028,n1029,n1030,n1031,n1032,n1033,n1034,n1035,
n1036,n1037,n1038,n1039,n1040,n1041,n1042,n1043,n1044,n1045,
n1046,n1047,n1048,n1049,n1050,n1051,n1052,n1053,n1054,n1055,
n1056,n1057,n1058,n1059,n1060,n1061,n1062,n1063,n1064,n1065,
n1066,n1067,n1068,n1069,n1070,n1071,n1072,n1073,n1074,n1075,
n1076,n1077,n1078,n1079,n1080,n1081,n1082,n1083,n1084,n1085,
n1086,n1087,n1088,n1089,n1090,n1091,n1092,n1093,n1094,n1095,
n1096,n1097,n1098,n1099,n1100,n1101,n1102,n1103,n1104,n1105,
n1106,n1107,n1108,n1109,n1110,n1111,n1112,n1113,n1114,n1115,
n1116,n1117,n1118,n1119,n1120,n1121,n1122,n1123,n1124,n1125,
n1126,n1127,n1128,n1129,n1130,n1131,n1132,n1133,n1134,n1135,
n1136,n1137,n1138,n1139,n1140,n1141,n1142,n1143,n1144,n1145,
n1146,n1147,n1148,n1149,n1150,n1151,n1152,n1153,n1154,n1155,
n1156,n1157,n1158,n1159,n1160,n1161,n1162,n1163,n1164,n1165,
n1166,n1167,n1168,n1169,n1170,n1171,n1172,n1173,n1174,n1175,
n1176,n1177,n1178,n1179,n1180,n1181,n1182,n1183,n1184,n1185,
n1186,n1187,n1188,n1189,n1190,n1191,n1192,n1193,n1194,n1195,
n1196,n1197,n1198,n1199,n1200,n1201,n1202,n1203,n1204,n1205,
n1206,n1207,n1208,n1210,n1211,n1212,n1213,n1214,n1216,n1217,
n1218,n1219,n1220,n1221,n1222,n1223,n1224,n1225,n1226,n1227,
n1228,n1229,n1230,n1231,n1232,n1233,n1234,n1235,n1236,n1237,
n1238,n1239,n1240,n1241,n1242,n1243,n1244,n1245,n1246,n1247,
n1248,n1249,n1250,n1251,n1252,n1253,n1254,n1255,n1256,n1257,
n1258,n1259,n1260,n1261,n1262,n1263,n1264,n1265,n1266,n1267,
n1268,n1269,n1270,n1271,n1272,n1273,n1274,n1275,n1276,n1277,
n1278,n1279,n1280,n1281,n1282,n1283,n1284,n1285,n1286,n1287,
n1288,n1289,n1290,n1291,n1292,n1293,n1294,n1295,n1296,n1297,
n1298,n1299,n1300,n1301,n1302,n1303,n1304,n1305,n1306,n1307,
n1308,n1309,n1310,n1311,n1312,n1313,n1314,n1315,n1316,n1317,
n1318,n1319,n1320,n1321,n1322,n1323,n1324,n1325,n1326,n1327,
n1328,n1329,n1330,n1331,n1332,n1333,n1334,n1335,n1336,n1337,
n1338,n1339,n1340,n1341,n1342,n1343,n1344,n1345,n1346,n1347,
n1348,n1349,n1350,n1351,n1352,n1353,n1354,n1355,n1356,n1357,
n1358,n1359,n1360,n1361,n1362,n1363,n1364,n1365,n1366,n1367,
n1368,n1369,n1370,n1371,n1372,n1373,n1374,n1375,n1376,n1377,
n1378,n1379,n1380,n1381,n1382,n1383,n1384,n1385,n1386,n1387,
n1388,n1389,n1390,n1391,n1392,n1393,n1394,n1395,n1396,n1397,
n1398,n1399,n1400,n1401,n1402,n1403,n1404,n1405,n1406,n1407,
n1408,n1409,n1410,n1411,n1412,n1413,n1414,n1415,n1416,n1417,
n1419,n1420,n1421,n1422,n1423,n1425,n1426,n1427,n1428,n1429,
n1430,n1431,n1432,n1433,n1434,n1435,n1436,n1437,n1438,n1439,
n1440,n1441,n1442,n1443,n1444,n1445,n1446,n1447,n1448,n1449,
n1450,n1451,n1452,n1453,n1454,n1455,n1456,n1457,n1458,n1459,
n1460,n1461,n1462,n1463,n1464,n1465,n1466,n1467,n1468,n1469,
n1470,n1471,n1472,n1473,n1474,n1475,n1476,n1477,n1478,n1479,
n1480,n1481,n1482,n1483,n1484,n1485,n1486,n1487,n1488,n1489,
n1490,n1491,n1492,n1493,n1494,n1495,n1496,n1497,n1498,n1499,
n1500,n1501,n1502,n1503,n1504,n1505,n1506,n1507,n1509,n1510,
n1511,n1512,n1513,n1515,n1516,n1517,n1518,n1519,n1520,n1521,
n1522,n1523,n1524,n1525,n1526,n1527,n1528,n1529,n1530,n1531,
n1532,n1533,n1534,n1535,n1536,n1537,n1538,n1539,n1540,n1541,
n1542,n1543,n1544,n1545,n1546,n1547,n1548,n1549,n1550,n1551,
n1552,n1553,n1554,n1555,n1556,n1557,n1558,n1559,n1560,n1561,
n1562,n1563,n1564,n1565,n1566,n1567,n1568,n1569,n1570,n1571,
n1572,n1573,n1574,n1575,n1576,n1577,n1578,n1579,n1580,n1581,
n1582,n1583,n1584,n1585,n1586,n1587,n1588,n1589,n1590,n1591,
n1592,n1593,n1594,n1595,n1596,n1597,n1598,n1599,n1600,n1601,
n1602,n1603,n1604,n1605,n1606,n1607,n1608,n1609,n1610,n1611,
n1612,n1613,n1614,n1615,n1616,n1617,n1618,n1619,n1620,n1621,
n1622,n1623,n1624,n1625,n1626,n1627,n1628,n1629,n1630,n1631,
n1632,n1633,n1634,n1635,n1636,n1637,n1638,n1639,n1640,n1641,
n1642,n1643,n1644,n1645,n1646,n1647,n1648,n1649,n1650,n1651,
n1652,n1653,n1654,n1655,n1656,n1657,n1658,n1659,n1660,n1661,
n1662,n1663,n1664,n1665,n1666,n1667,n1668,n1669,n1670,n1671,
n1672,n1673,n1674,n1675,n1676,n1677,n1678,n1679,n1680,n1681,
n1682,n1683,n1684,n1685,n1686,n1687,n1688,n1689,n1690,n1691,
n1692,n1693,n1694,n1695,n1696,n1697,n1698,n1699,n1700,n1701,
n1702,n1703,n1704,n1705,n1706,n1707,n1708,n1709,n1710,n1711,
n1712,n1713,n1715,n1716,n1717,n1718,n1719,n1721,n1722,n1723,
n1724,n1725,n1726,n1727,n1728,n1729,n1730,n1731,n1732,n1733,
n1734,n1735,n1736,n1737,n1738,n1739,n1740,n1741,n1742,n1743,
n1744,n1745,n1746,n1747,n1748,n1749,n1750,n1751,n1752,n1753,
n1754,n1755,n1756,n1757,n1758,n1759,n1760,n1761,n1762,n1763,
n1764,n1765,n1766,n1767,n1768,n1769,n1770,n1771,n1772,n1773,
n1774,n1775,n1776,n1777,n1778,n1779,n1780,n1781,n1782,n1783,
n1784,n1785,n1786,n1787,n1788,n1789,n1790,n1791,n1792,n1793,
n1794,n1795,n1796,n1797,n1798,n1799,n1800,n1801,n1802,n1803,
n1804,n1805,n1806,n1807,n1808,n1809,n1810,n1812,n1813,n1814,
n1815,n1816,n1817,n1818,n1819,n1820,n1821,n1822,n1824,n1825,
n1826,n1827,n1828,n1829,n1830,n1831,n1832,n1833,n1834,n1835,
n1836,n1837,n1838,n1839,n1840,n1841,n1842,n1843,n1844,n1845,
n1846,n1847,n1848,n1849,n1850,n1851,n1852,n1853,n1854,n1855,
n1856,n1857,n1858,n1859,n1860,n1861,n1862,n1863,n1864,n1865,
n1866,n1867,n1868,n1869,n1870,n1871,n1872,n1873,n1874,n1875,
n1876,n1877,n1878,n1879,n1880,n1881,n1882,n1883,n1884,n1885,
n1886,n1887,n1888,n1889,n1890,n1891,n1892,n1893,n1894,n1895,
n1896,n1897,n1898,n1899,n1900,n1901,n1902,n1903,n1904,n1905,
n1906,n1907,n1908,n1909,n1910,n1911,n1912,n1913,n1914,n1915,
n1916,n1917,n1918,n1919,n1920,n1921,n1922,n1923,n1924,n1925,
n1926,n1927,n1928,n1929,n1930,n1931,n1932,n1933,n1934,n1935,
n1936,n1937,n1938,n1939,n1940,n1941,n1942,n1943,n1944,n1945,
n1946,n1947,n1948,n1949,n1950,n1951,n1952,n1953,n1954,n1955,
n1956,n1957,n1958,n1959,n1960,n1961,n1962,n1963,n1964,n1965,
n1966,n1967,n1968,n1969,n1970,n1971,n1972,n1973,n1974,n1975,
n1976,n1977,n1978,n1979,n1980,n1981,n1982,n1983,n1984,n1985,
n1986,n1987,n1988,n1989,n1990,n1991,n1992,n1993,n1994,n1995,
n1996,n1997,n1998,n1999,n2000,n2001,n2002,n2003,n2004,n2005,
n2006,n2007,n2008,n2009,n2010,n2011,n2012,n2013,n2014,n2015,
n2016,n2017,n2018,n2019,n2020,n2021,n2022,n2023,n2024,n2025,
n2026,n2027,n2028,n2029,n2030,n2031,n2032,n2033,n2034,n2036,
n2037,n2038,n2039,n2040,n2041,n2042,n2043,n2044,n2045,n2046,
n2048,n2049,n2050,n2051,n2052,n2053,n2054,n2055,n2056,n2057,
n2058,n2059,n2060,n2061,n2062,n2063,n2064,n2065,n2066,n2067,
n2068,n2069,n2070,n2071,n2072,n2073,n2074,n2075,n2076,n2077,
n2078,n2079,n2080,n2081,n2082,n2083,n2084,n2085,n2086,n2087,
n2088,n2089,n2090,n2091,n2092,n2093,n2094,n2095,n2096,n2097,
n2098,n2099,n2100,n2101,n2102,n2103,n2104,n2105,n2106,n2107,
n2108,n2109,n2110,n2111,n2112,n2114,n2115,n2116,n2117,n2118,
n2119,n2120,n2121,n2122,n2123,n2124,n2126,n2127,n2128,n2129,
n2130,n2131,n2132,n2133,n2134,n2135,n2136,n2137,n2138,n2139,
n2140,n2141,n2142,n2143,n2144,n2145,n2146,n2147,n2148,n2149,
n2150,n2151,n2152,n2153,n2154,n2155,n2156,n2157,n2158,n2159,
n2160,n2161,n2162,n2163,n2164,n2165,n2166,n2167,n2168,n2169,
n2170,n2171,n2172,n2173,n2174,n2175,n2176,n2177,n2178,n2179,
n2180,n2181,n2182,n2183,n2184,n2185,n2186,n2187,n2188,n2189,
n2190,n2191,n2192,n2193,n2194,n2195,n2196,n2197,n2198,n2199,
n2200,n2201,n2202,n2203,n2204,n2205,n2206,n2207,n2208,n2209,
n2210,n2211,n2213,n2214,n2215,n2216,n2217,n2218,n2219,n2220,
n2221,n2222,n2223,n2225,n2226,n2227,n2228,n2229,n2230,n2231,
n2232,n2233,n2234,n2235,n2236,n2237,n2238,n2239,n2240,n2241,
n2242,n2243,n2244,n2245,n2246,n2247,n2248,n2249,n2250,n2251,
n2252,n2253,n2254,n2255,n2256,n2257,n2258,n2259,n2260,n2261,
n2262,n2263,n2264,n2265,n2266,n2267,n2268,n2269,n2270,n2271,
n2272,n2273,n2274,n2275,n2276,n2277,n2278,n2279,n2280,n2281,
n2282,n2283,n2284,n2285,n2286,n2287,n2288,n2289,n2290,n2291,
n2292,n2293,n2294,n2295,n2296,n2297,n2298,n2299,n2300,n2301,
n2302,n2303,n2304,n2305,n2306,n2307,n2308,n2309,n2310,n2311,
n2312,n2313,n2314,n2315,n2316,n2317,n2318,n2319,n2320,n2321,
n2322,n2323,n2324,n2325,n2326,n2327,n2328,n2329,n2330,n2331,
n2332,n2333,n2334,n2335,n2336,n2337,n2338,n2339,n2340,n2341,
n2342,n2343,n2344,n2345,n2346,n2347,n2348,n2349,n2350,n2351,
n2352,n2353,n2354,n2355,n2356,n2357,n2358,n2359,n2360,n2361,
n2362,n2363,n2364,n2365,n2366,n2367,n2368,n2369,n2370,n2371,
n2372,n2373,n2374,n2375,n2376,n2377,n2378,n2379,n2380,n2381,
n2382,n2383,n2384,n2385,n2386,n2387,n2388,n2389,n2390,n2391,
n2392,n2393,n2394,n2395,n2396,n2397,n2398,n2399,n2400,n2401,
n2402,n2403,n2404,n2405,n2406,n2407,n2408,n2409,n2410,n2411,
n2412,n2413,n2414,n2415,n2416,n2417,n2418,n2419,n2420,n2421,
n2422,n2423,n2424,n2425,n2426,n2427,n2428,n2429,n2430,n2431,
n2433,n2434,n2435,n2436,n2437,n2438,n2439,n2440,n2441,n2442,
n2443,n2445,n2446,n2447,n2448,n2449,n2450,n2451,n2452,n2453,
n2454,n2455,n2456,n2457,n2458,n2459,n2460,n2461,n2462,n2463,
n2464,n2465,n2466,n2467,n2468,n2469,n2470,n2471,n2472,n2473,
n2474,n2475,n2476,n2477,n2478,n2479,n2480,n2481,n2482,n2483,
n2484,n2485,n2486,n2487,n2488,n2489,n2490,n2491,n2492,n2493,
n2494,n2495,n2496,n2497,n2498,n2499,n2500,n2501,n2502,n2503,
n2504,n2505,n2506,n2507,n2508,n2509,n2510,n2511,n2512,n2513,
n2514,n2515,n2516,n2517,n2518,n2519,n2520,n2521,n2522,n2523,
n2524,n2525,n2526,n2527,n2528,n2529,n2530,n2531,n2532,n2533,
n2534,n2535,n2536,n2537,n2538,n2539,n2540,n2541,n2542,n2543,
n2544,n2545,n2546,n2547,n2548,n2549,n2550,n2551,n2552,n2553,
n2554,n2555,n2556,n2557,n2558,n2559,n2560,n2561,n2562,n2563,
n2564,n2565,n2566,n2567,n2568,n2569,n2570,n2571,n2572,n2573,
n2574,n2575,n2576,n2577,n2578,n2579,n2580,n2581,n2582,n2583,
n2584,n2585,n2586,n2587,n2588,n2589,n2590,n2591,n2592,n2593,
n2594,n2595,n2596,n2597,n2598,n2599,n2600,n2601,n2602,n2603,
n2604,n2605,n2606,n2607,n2608,n2609,n2610,n2611,n2612,n2613,
n2614,n2615,n2616,n2617,n2618,n2619,n2620,n2621,n2622,n2623,
n2624,n2625,n2626,n2627,n2628,n2629,n2630,n2631,n2632,n2633,
n2634,n2635,n2636,n2637,n2638,n2639,n2640,n2641,n2642,n2643,
n2644,n2645,n2646,n2647,n2648,n2650,n2651,n2652,n2653,n2654,
n2655,n2656,n2657,n2658,n2659,n2660,n2662,n2663,n2664,n2665,
n2666,n2667,n2668,n2669,n2670,n2671,n2672,n2673,n2674,n2675,
n2676,n2677,n2678,n2679,n2680,n2681,n2682,n2683,n2684,n2685,
n2686,n2687,n2688,n2689,n2690,n2691,n2692,n2693,n2694,n2695,
n2696,n2697,n2698,n2699,n2700,n2701,n2702,n2703,n2704,n2705,
n2706,n2707,n2708,n2709,n2710,n2711,n2712,n2713,n2714,n2715,
n2716,n2717,n2718,n2719,n2720,n2721,n2722,n2723,n2724,n2725,
n2726,n2727,n2728,n2729,n2730,n2731,n2732,n2733,n2734,n2735,
n2736,n2737,n2738,n2739,n2740,n2742,n2743,n2744,n2745,n2746,
n2747,n2748,n2749,n2750,n2751,n2752,n2754,n2755,n2756,n2757,
n2758,n2759,n2760,n2761,n2762,n2763,n2764,n2765,n2766,n2767,
n2768,n2769,n2770,n2771,n2772,n2773,n2774,n2775,n2776,n2777,
n2778,n2779,n2780,n2781,n2782,n2783,n2784,n2785,n2786,n2787,
n2788,n2789,n2790,n2791,n2792,n2793,n2794,n2795,n2796,n2797,
n2798,n2799,n2800,n2801,n2802,n2803,n2804,n2805,n2806,n2807,
n2808,n2809,n2810,n2811,n2812,n2813,n2814,n2815,n2816,n2817,
n2818,n2819,n2820,n2821,n2822,n2823,n2824,n2825,n2826,n2827,
n2828,n2829,n2830,n2831,n2832,n2833,n2834,n2835,n2836,n2837,
n2838,n2839,n2840,n2841,n2842,n2843,n2844,n2845,n2847,n2848,
n2849,n2850,n2851,n2852,n2853,n2854,n2855,n2856,n2857,n2859,
n2860,n2861,n2862,n2863,n2864,n2865,n2866,n2867,n2868,n2869,
n2870,n2871,n2872,n2873,n2874,n2875,n2876,n2877,n2878,n2879,
n2880,n2881,n2882,n2883,n2884,n2885,n2886,n2887,n2888,n2889,
n2890,n2891,n2892,n2893,n2894,n2895,n2896,n2897,n2898,n2899,
n2900,n2901,n2902,n2903,n2904,n2905,n2906,n2907,n2908,n2909,
n2910,n2911,n2912,n2913,n2915,n2916,n2917,n2918,n2919,n2920,
n2921,n2922,n2923,n2924,n2925,n2927,n2928,n2929,n2930,n2931,
n2932,n2933,n2934,n2935,n2936,n2937,n2938,n2939,n2940,n2941,
n2942,n2943,n2944,n2945,n2946,n2947,n2948,n2949,n2950,n2951,
n2952,n2953,n2954,n2955,n2956,n2957,n2958,n2959,n2960,n2961,
n2962,n2963,n2964,n2965,n2966,n2967,n2968,n2969,n2970,n2971,
n2972,n2973,n2974,n2975,n2976,n2977,n2978,n2980,n2981,n2982,
n2983,n2984,n2985,n2986,n2987,n2988,n2989,n2990,n2992,n2993,
n2994,n2995,n2996,n2997,n2998,n2999,n3000,n3001,n3002,n3003,
n3004,n3005,n3006,n3007,n3008,n3009,n3010,n3011,n3012,n3013,
n3014,n3015,n3016,n3017,n3018,n3019,n3020,n3021,n3022,n3023,
n3024,n3025,n3026,n3027,n3028,n3029,n3030,n3031,n3032,n3033,
n3034,n3035,n3036,n3037,n3038,n3039,n3040,n3041,n3042,n3043,
n3044,n3045,n3046,n3047,n3048,n3049,n3050,n3051,n3052,n3053,
n3054,n3055,n3056,n3057,n3058,n3059,n3060,n3061,n3062,n3063,
n3064,n3065,n3066,n3067,n3068,n3069,n3070,n3071,n3072,n3073,
n3074,n3075,n3076,n3077,n3078,n3079,n3080,n3081,n3082,n3083,
n3084,n3085,n3086,n3087,n3088,n3089,n3090,n3091,n3092,n3093,
n3094,n3095,n3096,n3097,n3098,n3099,n3100,n3101,n3102,n3103,
n3104,n3105,n3106,n3107,n3108,n3109,n3110,n3111,n3112,n3113,
n3114,n3115,n3116,n3117,n3118,n3119,n3120,n3121,n3122,n3123,
n3124,n3125,n3126,n3127,n3128,n3129,n3130,n3131,n3132,n3133,
n3134,n3135,n3136,n3137,n3138,n3139,n3140,n3141,n3142,n3143,
n3144,n3145,n3146,n3147,n3148,n3149,n3150,n3151,n3152,n3153,
n3154,n3155,n3156,n3157,n3158,n3159,n3160,n3161,n3162,n3163,
n3164,n3165,n3166,n3167,n3168,n3169,n3170,n3171,n3172,n3173,
n3174,n3175,n3176,n3177,n3178,n3179,n3180,n3181,n3182,n3183,
n3184,n3185,n3186,n3187,n3188,n3189,n3190,n3192,n3193,n3194,
n3195,n3196,n3197,n3198,n3199,n3200,n3201,n3202,n3204,n3205,
n3206,n3207,n3208,n3209,n3210,n3211,n3212,n3213,n3214,n3215,
n3216,n3217,n3218,n3219,n3220,n3221,n3222,n3223,n3224,n3225,
n3226,n3227,n3228,n3229,n3230,n3231,n3232,n3233,n3234,n3235,
n3236,n3237,n3238,n3239,n3240,n3241,n3242,n3243,n3244,n3245,
n3246,n3247,n3248,n3249,n3250,n3251,n3252,n3253,n3254,n3255,
n3256,n3257,n3258,n3259,n3260,n3261,n3262,n3263,n3264,n3265,
n3266,n3267,n3268,n3269,n3270,n3271,n3272,n3273,n3274,n3275,
n3276,n3277,n3279,n3280,n3281,n3282,n3283,n3284,n3285,n3286,
n3287,n3288,n3289,n3291,n3292,n3293,n3294,n3295,n3296,n3297,
n3298,n3299,n3300,n3301,n3302,n3303,n3304,n3305,n3306,n3307,
n3308,n3309,n3310,n3311,n3312,n3313,n3314,n3315,n3316,n3317,
n3318,n3319,n3320,n3321,n3322,n3323,n3324,n3325,n3326,n3327,
n3328,n3329,n3330,n3331,n3332,n3333,n3334,n3335,n3336,n3337,
n3338,n3339,n3340,n3341,n3342,n3343,n3344,n3346,n3347,n3348,
n3349,n3350,n3351,n3352,n3353,n3354,n3355,n3356,n3358,n3359,
n3360,n3361,n3362,n3363,n3364,n3365,n3366,n3367,n3368,n3369,
n3370,n3371,n3372,n3373,n3374,n3375,n3376,n3377,n3378,n3379,
n3380,n3381,n3382,n3383,n3384,n3385,n3386,n3387,n3388,n3389,
n3390,n3391,n3392,n3393,n3394,n3395,n3396,n3397,n3398,n3399,
n3400,n3401,n3402,n3403,n3404,n3405,n3406,n3407,n3408,n3409,
n3410,n3411,n3412,n3413,n3414,n3415,n3416,n3417,n3418,n3419,
n3420,n3421,n3422,n3423,n3424,n3425,n3426,n3427,n3428,n3429,
n3430,n3431,n3432,n3433,n3434,n3435,n3436,n3437,n3438,n3439,
n3440,n3441,n3442,n3443,n3444,n3445,n3447,n3448,n3449,n3450,
n3451,n3452,n3453,n3454,n3455,n3456,n3457,n3459,n3460,n3461,
n3462,n3463,n3464,n3465,n3466,n3467,n3468,n3469,n3470,n3471,
n3472,n3473,n3474,n3475,n3476,n3477,n3478,n3479,n3480,n3481,
n3482,n3483,n3484,n3485,n3486,n3487,n3488,n3489,n3490,n3491,
n3492,n3493,n3494,n3495,n3496,n3497,n3498,n3499,n3500,n3501,
n3502,n3503,n3504,n3505,n3506,n3507,n3508,n3509,n3510,n3511,
n3512,n3513,n3514,n3515,n3516,n3517,n3518,n3519,n3520,n3521,
n3522,n3523,n3524,n3525,n3526,n3527,n3529,n3530,n3531,n3532,
n3533,n3534,n3535,n3536,n3537,n3538,n3539,n3541,n3542,n3543,
n3544,n3545,n3546,n3547,n3548,n3549,n3550,n3551,n3552,n3553,
n3554,n3555,n3556,n3557,n3558,n3559,n3560,n3561,n3562,n3563,
n3564,n3565,n3566,n3567,n3568,n3569,n3570,n3571,n3572,n3573,
n3574,n3575,n3576,n3577,n3578,n3579,n3580,n3581,n3582,n3583,
n3584,n3585,n3586,n3587,n3588,n3589,n3590,n3591,n3592,n3593,
n3594,n3595,n3596,n3597,n3598,n3599,n3600,n3601,n3602,n3603,
n3605,n3606,n3607,n3608,n3609,n3610,n3611,n3612,n3613,n3614,
n3615,n3617,n3618,n3619,n3620,n3621,n3622,n3623,n3624,n3625,
n3626,n3627,n3628,n3629,n3630,n3631,n3632,n3633,n3634,n3635,
n3636,n3637,n3638,n3639,n3640,n3641,n3642,n3643,n3644,n3645,
n3646,n3647,n3648,n3649,n3650,n3651,n3652,n3653,n3654,n3655,
n3656,n3657,n3658,n3659,n3660,n3661,n3662,n3663,n3664,n3665,
n3666,n3667,n3668,n3669,n3670,n3671,n3672,n3673,n3674,n3675,
n3676,n3677,n3678,n3679,n3680,n3681,n3682,n3683,n3684,n3685,
n3686,n3687,n3688,n3689,n3690,n3691,n3692,n3693,n3694,n3695,
n3696,n3697,n3698,n3699,n3700,n3701,n3702,n3703,n3704,n3705,
n3706,n3707,n3708,n3709,n3710,n3711,n3712,n3713,n3714,n3715,
n3716,n3717,n3718,n3719,n3720,n3721,n3722,n3723,n3724,n3725,
n3726,n3727,n3728,n3729,n3730,n3731,n3732,n3733,n3734,n3735,
n3736,n3737,n3738,n3739,n3740,n3741,n3742,n3743,n3744,n3745,
n3746,n3747,n3748,n3749,n3750,n3751,n3752,n3753,n3754,n3755,
n3756,n3757,n3758,n3759,n3760,n3761,n3762,n3763,n3764,n3765,
n3766,n3767,n3768,n3769,n3770,n3771,n3772,n3773,n3774,n3775,
n3776,n3777,n3778,n3779,n3780,n3781,n3782,n3783,n3784,n3785,
n3786,n3787,n3788,n3789,n3790,n3791,n3792,n3793,n3794,n3795,
n3796,n3797,n3798,n3799,n3800,n3801,n3802,n3803,n3804,n3805,
n3806,n3807,n3808,n3809,n3810,n3811,n3812,n3813,n3814,n3815,
n3816,n3817,n3818,n3819,n3820,n3821,n3822,n3824,n3825,n3826,
n3827,n3828,n3829,n3830,n3831,n3832,n3833,n3834,n3836,n3837,
n3838,n3839,n3840,n3841,n3842,n3843,n3844,n3845,n3846,n3847,
n3848,n3849,n3850,n3851,n3852,n3853,n3854,n3855,n3856,n3857,
n3858,n3859,n3860,n3861,n3862,n3863,n3864,n3865,n3866,n3867,
n3868,n3869,n3870,n3871,n3872,n3873,n3874,n3875,n3876,n3877,
n3878,n3879,n3880,n3881,n3882,n3883,n3884,n3885,n3886,n3887,
n3888,n3889,n3890,n3891,n3892,n3893,n3894,n3895,n3896,n3897,
n3898,n3899,n3900,n3901,n3902,n3903,n3904,n3905,n3906,n3907,
n3908,n3909,n3910,n3911,n3912,n3913,n3914,n3915,n3916,n3917,
n3918,n3919,n3920,n3922,n3923,n3924,n3925,n3926,n3927,n3928,
n3929,n3930,n3931,n3932,n3934,n3935,n3936,n3937,n3938,n3939,
n3940,n3941,n3942,n3943,n3944,n3945,n3946,n3947,n3948,n3949,
n3950,n3951,n3952,n3953,n3954,n3955,n3956,n3957,n3958,n3959,
n3960,n3961,n3962,n3963,n3964,n3965,n3966,n3967,n3968,n3969,
n3970,n3971,n3972,n3973,n3974,n3975,n3976,n3977,n3978,n3979,
n3980,n3981,n3982,n3983,n3984,n3985,n3986,n3987,n3988,n3989,
n3990,n3991,n3992,n3993,n3994,n3995,n3996,n3997,n3998,n3999,
n4000,n4001,n4002,n4003,n4004,n4006,n4007,n4008,n4009,n4010,
n4011,n4012,n4013,n4014,n4015,n4016,n4018,n4019,n4020,n4021,
n4022,n4023,n4024,n4025,n4026,n4027,n4028,n4029,n4030,n4031,
n4032,n4033,n4034,n4035,n4036,n4037,n4038,n4039,n4040,n4041,
n4042,n4043,n4044,n4045,n4046,n4047,n4048,n4049,n4050,n4051,
n4052,n4053,n4054,n4055,n4056,n4057,n4058,n4059,n4060,n4061,
n4062,n4063,n4064,n4065,n4066,n4067,n4068,n4069,n4070,n4071,
n4072,n4073,n4074,n4075,n4076,n4077,n4078,n4079,n4080,n4081,
n4082,n4083,n4084,n4085,n4086,n4087,n4088,n4089,n4090,n4091,
n4092,n4093,n4094,n4095,n4096,n4097,n4098,n4099,n4100,n4101,
n4102,n4103,n4104,n4105,n4106,n4108,n4109,n4110,n4111,n4112,
n4113,n4114,n4115,n4116,n4117,n4118,n4120,n4121,n4122,n4123,
n4124,n4125,n4126,n4127,n4128,n4129,n4130,n4131,n4132,n4133,
n4134,n4135,n4136,n4137,n4138,n4139,n4140,n4141,n4142,n4143,
n4144,n4145,n4146,n4147,n4148,n4149,n4150,n4151,n4152,n4153,
n4154,n4155,n4156,n4157,n4158,n4159,n4160,n4161,n4162,n4163,
n4164,n4165,n4166,n4167,n4168,n4169,n4170,n4171,n4172,n4173,
n4174,n4175,n4176,n4177,n4178,n4179,n4180,n4181,n4182,n4183,
n4184,n4185,n4186,n4187,n4189,n4190,n4191,n4192,n4193,n4194,
n4195,n4196,n4197,n4198,n4199,n4201,n4202,n4203,n4204,n4205,
n4206,n4207,n4208,n4209,n4210,n4211,n4212,n4213,n4214,n4215,
n4216,n4217,n4218,n4219,n4220,n4221,n4222,n4223,n4224,n4225,
n4226,n4227,n4228,n4229,n4230,n4231,n4232,n4233,n4234,n4235,
n4236,n4237,n4238,n4239,n4240,n4241,n4242,n4243,n4244,n4245,
n4246,n4247,n4248,n4249,n4250,n4251,n4253,n4254,n4255,n4256,
n4257,n4258,n4259,n4260,n4261,n4262,n4263,n4265,n4266,n4267,
n4268,n4269,n4270,n4271,n4272,n4273,n4274,n4275,n4276,n4277,
n4278,n4279,n4280,n4281,n4282,n4283,n4284,n4285,n4286,n4287,
n4288,n4289,n4290,n4291,n4292,n4293,n4294,n4295,n4296,n4297,
n4298,n4299,n4300,n4301,n4302,n4303,n4304,n4305,n4306,n4307,
n4308,n4309,n4310,n4311,n4312,n4313,n4314,n4315,n4316,n4317,
n4318,n4319,n4320,n4321,n4322,n4323,n4324,n4326,n4327,n4328,
n4329,n4330,n4331,n4332,n4333,n4334,n4335,n4336,n4338,n4339,
n4340,n4341,n4342,n4343,n4344,n4345,n4346,n4347,n4348,n4349,
n4350,n4351,n4352,n4353,n4354,n4355,n4356,n4357,n4358,n4359,
n4360,n4361,n4362,n4363,n4364,n4365,n4366,n4367,n4368,n4369,
n4370,n4371,n4372,n4373,n4374,n4375,n4376,n4377,n4378,n4379,
n4380,n4381,n4382,n4383,n4384,n4385,n4386,n4387,n4388,n4389,
n4390,n4391,n4392,n4393,n4394,n4395,n4396,n4397,n4398,n4399,
n4400,n4401,n4402,n4403,n4404,n4406,n4407,n4408,n4409,n4410,
n4411,n4412,n4413,n4414,n4415,n4416,n4418,n4419,n4420,n4421,
n4422,n4423,n4424,n4425,n4426,n4427,n4428,n4429,n4430,n4431,
n4432,n4433,n4434,n4435,n4436,n4437,n4438,n4439,n4440,n4441,
n4442,n4443,n4444,n4445,n4446,n4447,n4448,n4449,n4450,n4451,
n4452,n4453,n4454,n4455,n4456,n4457,n4458,n4459,n4460,n4461,
n4462,n4463,n4464,n4465,n4466,n4467,n4468,n4469,n4470,n4471,
n4472,n4473,n4474,n4475,n4477,n4478,n4479,n4480,n4481,n4482,
n4483,n4484,n4485,n4486,n4487,n4489,n4490,n4491,n4492,n4493,
n4494,n4495,n4496,n4497,n4498,n4499,n4500,n4501,n4502,n4503,
n4504,n4505,n4506,n4507,n4508,n4509,n4510,n4511,n4512,n4513,
n4514,n4515,n4516,n4517,n4518,n4519,n4520,n4521,n4522,n4523,
n4524,n4525,n4526,n4527,n4528,n4529,n4530,n4531,n4532,n4533,
n4534,n4535,n4536,n4537,n4538,n4539,n4540,n4541,n4542,n4543,
n4544,n4545,n4546,n4547,n4548,n4549,n4550,n4551,n4552,n4553,
n4554,n4556,n4557,n4558,n4559,n4560,n4561,n4562,n4563,n4564,
n4565,n4566,n4568,n4569,n4570,n4571,n4572,n4573,n4574,n4575,
n4576,n4577,n4578,n4579,n4580,n4581,n4582,n4583,n4584,n4585,
n4586,n4587,n4588,n4589,n4590,n4591,n4592,n4593,n4594,n4595,
n4596,n4597,n4598,n4599,n4600,n4601,n4602,n4603,n4604,n4605,
n4606,n4607,n4608,n4609,n4610,n4611,n4612,n4613,n4614,n4615,
n4617,n4618,n4619,n4620,n4621,n4622,n4623,n4624,n4625,n4626,
n4627,n4629,n4630,n4631,n4632,n4633,n4634,n4635,n4636,n4637,
n4638,n4639,n4640,n4641,n4642,n4643,n4644,n4645,n4646,n4647,
n4648,n4649,n4650,n4651,n4652,n4653,n4654,n4655,n4656,n4657,
n4658,n4659,n4660,n4661,n4662,n4663,n4664,n4665,n4666,n4667,
n4668,n4669,n4670,n4671,n4672,n4673,n4674,n4675,n4676,n4677,
n4678,n4679,n4680,n4682,n4683,n4684,n4685,n4686,n4687,n4688,
n4689,n4690,n4691,n4692,n4694,n4695,n4696,n4697,n4698,n4700,
n4701,n4702,n4703,n4704,n4706,n4707,n4708,n4709,n4710,n4712,
n4713,n4714,n4715,n4716,n4718,n4719,n4720,n4721,n4722,n4724,
n4725,n4726,n4727,n4728,n4730,n4731,n4732,n4733,n4734,n4736,
n4737,n4738,n4739,n4740,n4742,n4743,n4744,n4745,n4746,n4748,
n4749,n4750,n4751,n4752,n4754,n4755,n4756,n4757,n4758,n4760,
n4761,n4762,n4763,n4764,n4766,n4767,n4768,n4769,n4770,n4772,
n4773,n4774,n4775,n4776,n4778,n4779,n4780,n4781,n4782,n4784,
n4785,n4786,n4787,n4788,n4790,n4791,n4792,n4793,n4794,n4796,
n4797,n4798,n4799,n4800,n4802,n4803,n4804,n4805,n4806,n4808,
n4809,n4810,n4811,n4812,n4814,n4815,n4816,n4817,n4818,n4820,
n4821,n4822,n4823,n4824,n4826,n4827,n4828,n4829,n4830,n4832,
n4833,n4834,n4835,n4836,n4838,n4839,n4840,n4841,n4842,n4844,
n4845,n4846,n4847,n4848,n4850,n4851,n4852,n4853,n4854,n4856,
n4857,n4858,n4859,n4860,n4862,n4863,n4864,n4865,n4866,n4868,
n4869,n4870,n4871,n4872,n4874,n4875,n4876,n4877,n4878,n4880,
n4881,n4882,n4883,n4884,n4886,n4887,n4888,n4889,n4890,n4892,
n4893,n4894,n4895,n4896,n4898,n4899,n4900,n4901,n4902,n4904,
n4905,n4906,n4907,n4908,n4910,n4911,n4912,n4913,n4914,n4916,
n4917,n4918,n4919,n4920,n4922,n4923,n4924,n4925,n4926,n4928,
n4929,n4930,n4931,n4932,n4934,n4935,n4936,n4937,n4938,n4940,
n4941,n4942,n4943,n4944,n4946,n4947,n4948,n4949,n4950,n4952,
n4953,n4954,n4955,n4956,n4958,n4959,n4960,n4961,n4962,n4964,
n4965,n4966,n4967,n4968,n4970,n4971,n4972,n4973,n4974,n4976,
n4977,n4978,n4979,n4980,n4982,n4983,n4984,n4985,n4986,n4988,
n4989,n4990,n4991,n4992,n4994,n4995,n4996,n4997,n4998,n5000,
n5001,n5002,n5003,n5004,n5006,n5007,n5008,n5009,n5010,n5012,
n5013,n5014,n5015,n5016,n5018,n5019,n5020,n5021,n5022,n5024,
n5025,n5026,n5027,n5028,n5030,n5031,n5032,n5033,n5034,n5036,
n5037,n5038,n5039,n5040,n5042,n5043,n5044,n5045,n5046,n5048,
n5049,n5050,n5051,n5052,n5054,n5055,n5056,n5057,n5058,n5060,
n5061,n5062,n5063,n5064,n5066,n5067,n5068,n5069,n5070,n5072,
n5073,n5074,n5075,n5076,n5078,n5079,n5080,n5081,n5082,n5083,
n5084,n5085,n5086,n5087,n5088,n5090,n5091,n5092,n5094,n5095,
n5096,n5097,n5098,n5099,n5102,n5103,n5104,n5105,n5106,n5107,
n5108,n5109,n5110,n5111,n5112,n5113,n5114,n5115,n5116,n5117,
n5118,n5119,n5120,n5121,n5122,n5123,n5124,n5125,n5126,n5127,
n5128,n5129,n5130,n5131,n5132,n5133,n5134,n5135,n5136,n5137,
n5138,n5139,n5140,n5141,n5142,n5143,n5144,n5145,n5146,n5147,
n5148,n5149,n5150,n5151,n5152,n5153,n5154,n5155,n5157,n5158,
n5159,n5160,n5161,n5162,n5163,n5164,n5165,n5166,n5167,n5168,
n5169,n5170,n5171,n5172,n5173,n5174,n5175,n5176,n5177,n5178,
n5179,n5180,n5181,n5182,n5183,n5184,n5185,n5186,n5187,n5188,
n5189,n5190,n5191,n5192,n5194,n5195,n5196,n5197,n5198,n5199,
n5200,n5201,n5202,n5203,n5204,n5205,n5206,n5207,n5208,n5209,
n5210,n5211,n5212,n5213,n5214,n5215,n5216,n5217,n5218,n5219,
n5220,n5221,n5222,n5223,n5224,n5225,n5226,n5227,n5229,n5230,
n5231,n5232,n5233,n5234,n5235,n5236,n5237,n5238,n5239,n5240,
n5241,n5242,n5243,n5244,n5245,n5246,n5247,n5248,n5249,n5250,
n5251,n5252,n5253,n5254,n5255,n5256,n5257,n5258,n5259,n5260,
n5261,n5262,n5264,n5265,n5266,n5267,n5268,n5269,n5270,n5271,
n5272,n5273,n5274,n5275,n5276,n5277,n5278,n5279,n5280,n5281,
n5282,n5283,n5284,n5285,n5286,n5287,n5288,n5289,n5290,n5291,
n5292,n5293,n5294,n5295,n5297,n5298,n5299,n5300,n5301,n5302,
n5303,n5304,n5305,n5306,n5307,n5308,n5309,n5310,n5311,n5312,
n5313,n5314,n5315,n5316,n5317,n5318,n5319,n5320,n5321,n5322,
n5323,n5324,n5325,n5326,n5327,n5328,n5330,n5331,n5332,n5333,
n5334,n5335,n5336,n5337,n5338,n5339,n5340,n5341,n5342,n5343,
n5344,n5345,n5346,n5347,n5348,n5349,n5350,n5351,n5352,n5353,
n5354,n5355,n5356,n5357,n5358,n5359,n5360,n5361,n5363,n5364,
n5365,n5366,n5367,n5368,n5369,n5370,n5371,n5372,n5373,n5374,
n5375,n5376,n5377,n5378,n5379,n5380,n5381,n5382,n5383,n5384,
n5385,n5386,n5387,n5388,n5389,n5390,n5391,n5392,n5393,n5394,
n5396,n5397,n5398,n5399,n5400,n5401,n5402,n5403,n5404,n5405,
n5406,n5407,n5408,n5409,n5410,n5411,n5412,n5413,n5414,n5415,
n5416,n5417,n5418,n5419,n5420,n5421,n5422,n5423,n5424,n5425,
n5426,n5427,n5429,n5430,n5431,n5432,n5433,n5434,n5435,n5436,
n5437,n5438,n5439,n5440,n5441,n5442,n5443,n5444,n5445,n5446,
n5447,n5448,n5449,n5450,n5451,n5452,n5453,n5454,n5455,n5456,
n5457,n5458,n5459,n5460,n5462,n5463,n5464,n5465,n5466,n5467,
n5468,n5469,n5470,n5471,n5472,n5473,n5474,n5475,n5476,n5477,
n5478,n5479,n5480,n5481,n5482,n5483,n5484,n5485,n5486,n5487,
n5488,n5489,n5490,n5491,n5492,n5493,n5495,n5496,n5497,n5498,
n5499,n5500,n5501,n5502,n5503,n5504,n5505,n5506,n5507,n5508,
n5509,n5510,n5511,n5512,n5513,n5514,n5515,n5516,n5517,n5518,
n5519,n5520,n5521,n5522,n5523,n5524,n5525,n5526,n5528,n5529,
n5530,n5531,n5532,n5533,n5534,n5535,n5536,n5537,n5538,n5539,
n5540,n5541,n5542,n5543,n5544,n5545,n5546,n5547,n5548,n5549,
n5550,n5551,n5552,n5553,n5554,n5555,n5556,n5557,n5558,n5559,
n5561,n5562,n5563,n5564,n5565,n5566,n5567,n5568,n5569,n5570,
n5571,n5572,n5573,n5574,n5575,n5576,n5577,n5578,n5579,n5580,
n5581,n5582,n5583,n5584,n5585,n5586,n5587,n5588,n5589,n5590,
n5591,n5592,n5594,n5595,n5596,n5597,n5598,n5599,n5600,n5601,
n5602,n5603,n5604,n5605,n5606,n5607,n5608,n5609,n5610,n5611,
n5612,n5613,n5614,n5615,n5616,n5617,n5618,n5619,n5620,n5621,
n5622,n5623,n5624,n5625,n5627,n5628,n5629,n5630,n5631,n5632,
n5633,n5634,n5635,n5636,n5637,n5638,n5639,n5640,n5641,n5642,
n5643,n5644,n5645,n5646,n5647,n5648,n5649,n5650,n5651,n5652,
n5653,n5654,n5655,n5656,n5657,n5658,n5660,n5661,n5662,n5663,
n5664,n5665,n5666,n5667,n5668,n5669,n5670,n5671,n5672,n5673,
n5674,n5675,n5676,n5677,n5678,n5679,n5680,n5681,n5682,n5683,
n5684,n5685,n5686,n5687,n5688,n5689,n5690,n5691,n5693,n5694,
n5695,n5696,n5697,n5698,n5699,n5700,n5701,n5702,n5703,n5704,
n5705,n5706,n5707,n5708,n5709,n5710,n5711,n5712,n5713,n5714,
n5715,n5716,n5717,n5718,n5719,n5720,n5721,n5722,n5723,n5724,
n5726,n5727,n5728,n5729,n5730,n5731,n5732,n5733,n5734,n5735,
n5736,n5737,n5738,n5739,n5740,n5741,n5742,n5743,n5744,n5745,
n5746,n5747,n5748,n5749,n5750,n5751,n5752,n5753,n5754,n5755,
n5756,n5757,n5759,n5760,n5761,n5762,n5763,n5764,n5765,n5766,
n5767,n5768,n5769,n5770,n5771,n5772,n5773,n5774,n5775,n5776,
n5777,n5778,n5779,n5780,n5781,n5782,n5783,n5784,n5785,n5786,
n5787,n5788,n5789,n5790,n5792,n5793,n5794,n5795,n5796,n5797,
n5798,n5799,n5800,n5801,n5802,n5803,n5804,n5805,n5806,n5807,
n5808,n5809,n5810,n5811,n5812,n5813,n5814,n5815,n5816,n5817,
n5818,n5819,n5820,n5821,n5822,n5823,n5825,n5826,n5827,n5828,
n5829,n5830,n5831,n5832,n5833,n5834,n5835,n5836,n5837,n5838,
n5839,n5840,n5841,n5842,n5843,n5844,n5845,n5846,n5847,n5848,
n5849,n5850,n5851,n5852,n5853,n5854,n5855,n5856,n5858,n5859,
n5860,n5861,n5862,n5863,n5864,n5865,n5866,n5867,n5868,n5869,
n5870,n5871,n5872,n5873,n5874,n5875,n5876,n5877,n5878,n5879,
n5880,n5881,n5882,n5883,n5884,n5885,n5886,n5887,n5888,n5889,
n5891,n5892,n5893,n5894,n5895,n5896,n5897,n5898,n5899,n5900,
n5901,n5902,n5903,n5904,n5905,n5906,n5907,n5908,n5909,n5910,
n5911,n5912,n5913,n5914,n5915,n5916,n5917,n5918,n5919,n5920,
n5921,n5922,n5924,n5925,n5926,n5927,n5928,n5929,n5930,n5931,
n5932,n5933,n5934,n5935,n5936,n5937,n5938,n5939,n5940,n5941,
n5942,n5943,n5944,n5945,n5946,n5947,n5948,n5949,n5950,n5951,
n5952,n5953,n5955,n5956,n5957,n5958,n5959,n5960,n5961,n5962,
n5963,n5964,n5965,n5966,n5967,n5968,n5969,n5970,n5971,n5972,
n5973,n5974,n5975,n5976,n5977,n5978,n5979,n5980,n5981,n5982,
n5983,n5984,n5986,n5987,n5988,n5989,n5990,n5991,n5992,n5993,
n5994,n5995,n5996,n5997,n5998,n5999,n6000,n6001,n6002,n6003,
n6004,n6005,n6006,n6007,n6008,n6009,n6010,n6011,n6012,n6013,
n6015,n6016,n6017,n6018,n6019,n6020,n6021,n6022,n6023,n6024,
n6025,n6026,n6027,n6028,n6029,n6030,n6031,n6032,n6033,n6034,
n6035,n6036,n6037,n6038,n6039,n6040,n6041,n6042,n6044,n6045,
n6046,n6047,n6048,n6049,n6050,n6051,n6052,n6053,n6054,n6055,
n6056,n6057,n6058,n6059,n6060,n6061,n6062,n6063,n6064,n6065,
n6066,n6067,n6068,n6069,n6070,n6071,n6072,n6073,n6074,n6075,
n6076,n6077,n6078,n6079,n6081,n6082,n6083,n6084,n6085,n6086,
n6087,n6088,n6089,n6090,n6091,n6092,n6093,n6094,n6095,n6096,
n6097,n6098,n6099,n6100,n6101,n6102,n6103,n6104,n6105,n6106,
n6107,n6108,n6109,n6110,n6111,n6112,n6113,n6114,n6115,n6116,
n6118,n6119,n6120,n6121,n6122,n6123,n6124,n6125,n6126,n6127,
n6128,n6129,n6130,n6131,n6132,n6133,n6134,n6135,n6136,n6137,
n6138,n6139,n6140,n6141,n6142,n6143,n6144,n6145,n6146,n6147,
n6148,n6149,n6150,n6151,n6153,n6154,n6155,n6156,n6157,n6158,
n6159,n6160,n6161,n6162,n6163,n6164,n6165,n6166,n6167,n6168,
n6169,n6170,n6171,n6172,n6173,n6174,n6175,n6176,n6177,n6178,
n6179,n6180,n6181,n6182,n6183,n6184,n6185,n6186,n6188,n6189,
n6190,n6191,n6192,n6193,n6194,n6195,n6196,n6197,n6198,n6199,
n6200,n6201,n6202,n6203,n6204,n6205,n6206,n6207,n6208,n6209,
n6210,n6211,n6212,n6213,n6214,n6215,n6216,n6217,n6218,n6219,
n6221,n6222,n6223,n6224,n6225,n6226,n6227,n6228,n6229,n6230,
n6231,n6232,n6233,n6234,n6235,n6236,n6237,n6238,n6239,n6240,
n6241,n6242,n6243,n6244,n6245,n6246,n6247,n6248,n6249,n6250,
n6251,n6252,n6254,n6255,n6256,n6257,n6258,n6259,n6260,n6261,
n6262,n6263,n6264,n6265,n6266,n6267,n6268,n6269,n6270,n6271,
n6272,n6273,n6274,n6275,n6276,n6277,n6278,n6279,n6280,n6281,
n6282,n6283,n6284,n6285,n6287,n6288,n6289,n6290,n6291,n6292,
n6293,n6294,n6295,n6296,n6297,n6298,n6299,n6300,n6301,n6302,
n6303,n6304,n6305,n6306,n6307,n6308,n6309,n6310,n6311,n6312,
n6313,n6314,n6315,n6316,n6317,n6318,n6320,n6321,n6322,n6323,
n6324,n6325,n6326,n6327,n6328,n6329,n6330,n6331,n6332,n6333,
n6334,n6335,n6336,n6337,n6338,n6339,n6340,n6341,n6342,n6343,
n6344,n6345,n6346,n6347,n6348,n6349,n6350,n6351,n6353,n6354,
n6355,n6356,n6357,n6358,n6359,n6360,n6361,n6362,n6363,n6364,
n6365,n6366,n6367,n6368,n6369,n6370,n6371,n6372,n6373,n6374,
n6375,n6376,n6377,n6378,n6379,n6380,n6381,n6382,n6383,n6384,
n6386,n6387,n6388,n6389,n6390,n6391,n6392,n6393,n6394,n6395,
n6396,n6397,n6398,n6399,n6400,n6401,n6402,n6403,n6404,n6405,
n6406,n6407,n6408,n6409,n6410,n6411,n6412,n6413,n6414,n6415,
n6416,n6417,n6419,n6420,n6421,n6422,n6423,n6424,n6425,n6426,
n6427,n6428,n6429,n6430,n6431,n6432,n6433,n6434,n6435,n6436,
n6437,n6438,n6439,n6440,n6441,n6442,n6443,n6444,n6445,n6446,
n6447,n6448,n6449,n6450,n6452,n6453,n6454,n6455,n6456,n6457,
n6458,n6459,n6460,n6461,n6462,n6463,n6464,n6465,n6466,n6467,
n6468,n6469,n6470,n6471,n6472,n6473,n6474,n6475,n6476,n6477,
n6478,n6479,n6480,n6481,n6482,n6483,n6485,n6486,n6487,n6488,
n6489,n6490,n6491,n6492,n6493,n6494,n6495,n6496,n6497,n6498,
n6499,n6500,n6501,n6502,n6503,n6504,n6505,n6506,n6507,n6508,
n6509,n6510,n6511,n6512,n6513,n6514,n6515,n6516,n6518,n6519,
n6520,n6521,n6522,n6523,n6524,n6525,n6526,n6527,n6528,n6529,
n6530,n6531,n6532,n6533,n6534,n6535,n6536,n6537,n6538,n6539,
n6540,n6541,n6542,n6543,n6544,n6545,n6546,n6547,n6548,n6549,
n6551,n6552,n6553,n6554,n6555,n6556,n6557,n6558,n6559,n6560,
n6561,n6562,n6563,n6564,n6565,n6566,n6567,n6568,n6569,n6570,
n6571,n6572,n6573,n6574,n6575,n6576,n6577,n6578,n6579,n6580,
n6581,n6582,n6584,n6585,n6586,n6587,n6588,n6589,n6590,n6591,
n6592,n6593,n6594,n6595,n6596,n6597,n6598,n6599,n6600,n6601,
n6602,n6603,n6604,n6605,n6606,n6607,n6608,n6609,n6610,n6611,
n6612,n6613,n6614,n6615,n6617,n6618,n6619,n6620,n6621,n6622,
n6623,n6624,n6625,n6626,n6627,n6628,n6629,n6630,n6631,n6632,
n6633,n6634,n6635,n6636,n6637,n6638,n6639,n6640,n6641,n6642,
n6643,n6644,n6645,n6646,n6647,n6648,n6650,n6651,n6652,n6653,
n6654,n6655,n6656,n6657,n6658,n6659,n6660,n6661,n6662,n6663,
n6664,n6665,n6666,n6667,n6668,n6669,n6670,n6671,n6672,n6673,
n6674,n6675,n6676,n6677,n6678,n6679,n6680,n6681,n6683,n6684,
n6685,n6686,n6687,n6688,n6689,n6690,n6691,n6692,n6693,n6694,
n6695,n6696,n6697,n6698,n6699,n6700,n6701,n6702,n6703,n6704,
n6705,n6706,n6707,n6708,n6709,n6710,n6711,n6712,n6713,n6714,
n6716,n6717,n6718,n6719,n6720,n6721,n6722,n6723,n6724,n6725,
n6726,n6727,n6728,n6729,n6730,n6731,n6732,n6733,n6734,n6735,
n6736,n6737,n6738,n6739,n6740,n6741,n6742,n6743,n6744,n6745,
n6746,n6747,n6749,n6750,n6751,n6752,n6753,n6754,n6755,n6756,
n6757,n6758,n6759,n6760,n6761,n6762,n6763,n6764,n6765,n6766,
n6767,n6768,n6769,n6770,n6771,n6772,n6773,n6774,n6775,n6776,
n6777,n6778,n6779,n6780,n6782,n6783,n6784,n6785,n6786,n6787,
n6788,n6789,n6790,n6791,n6792,n6793,n6794,n6795,n6796,n6797,
n6798,n6799,n6800,n6801,n6802,n6803,n6804,n6805,n6806,n6807,
n6808,n6809,n6810,n6811,n6812,n6813,n6815,n6816,n6817,n6818,
n6819,n6820,n6821,n6822,n6823,n6824,n6825,n6826,n6827,n6828,
n6829,n6830,n6831,n6832,n6833,n6834,n6835,n6836,n6837,n6838,
n6839,n6840,n6841,n6842,n6843,n6844,n6845,n6846,n6848,n6849,
n6850,n6851,n6852,n6853,n6854,n6855,n6856,n6857,n6858,n6859,
n6860,n6861,n6862,n6863,n6864,n6865,n6866,n6867,n6868,n6869,
n6870,n6871,n6872,n6873,n6874,n6875,n6876,n6877,n6879,n6880,
n6881,n6882,n6883,n6884,n6885,n6886,n6887,n6888,n6889,n6890,
n6891,n6892,n6893,n6894,n6895,n6896,n6897,n6898,n6899,n6900,
n6901,n6902,n6903,n6904,n6905,n6906,n6907,n6908,n6910,n6911,
n6912,n6913,n6914,n6915,n6916,n6917,n6918,n6919,n6920,n6921,
n6922,n6923,n6924,n6925,n6926,n6927,n6928,n6929,n6930,n6931,
n6932,n6933,n6934,n6935,n6936,n6937,n6939,n6940,n6941,n6942,
n6943,n6944,n6945,n6946,n6947,n6948,n6949,n6950,n6951,n6952,
n6953,n6954,n6955,n6956,n6957,n6958,n6959,n6960,n6961,n6962,
n6963,n6964,n6965,n6966,n6968,n6969,n6970,n6971,n6972;
not gate_0(n501,pi008);
not gate_1(n502,pi009);
not gate_2(n503,pi131);
not gate_3(n504,pi132);
not gate_4(n505,pi133);
not gate_5(n506,pi134);
not gate_6(n507,pi135);
not gate_7(n508,pi136);
not gate_8(n509,pi137);
not gate_9(n510,pi138);
not gate_10(n511,pi139);
not gate_11(n512,pi140);
not gate_12(n513,pi141);
not gate_13(n514,pi142);
not gate_14(n515,pi143);
not gate_15(n516,pi144);
not gate_16(n517,pi145);
not gate_17(n518,pi146);
not gate_18(n519,pi147);
not gate_19(n520,pi148);
not gate_20(n521,pi149);
not gate_21(n522,pi150);
not gate_22(n523,pi151);
not gate_23(n524,pi152);
not gate_24(n525,pi153);
not gate_25(n526,pi154);
not gate_26(n527,pi155);
not gate_27(n528,pi156);
not gate_28(n529,pi157);
not gate_29(n530,pi158);
not gate_30(n531,pi159);
not gate_31(n532,pi160);
not gate_32(n533,pi161);
not gate_33(n534,pi162);
not gate_34(n535,pi163);
not gate_35(n536,pi164);
not gate_36(n537,pi165);
not gate_37(n538,pi166);
not gate_38(n539,pi167);
not gate_39(n540,pi168);
not gate_40(n541,pi169);
not gate_41(n542,pi170);
not gate_42(n543,pi171);
not gate_43(n544,pi172);
not gate_44(n545,pi173);
not gate_45(n546,pi174);
not gate_46(n547,pi175);
not gate_47(n548,pi176);
not gate_48(n549,pi177);
not gate_49(n550,pi178);
not gate_50(n551,pi179);
not gate_51(n552,pi180);
not gate_52(n553,pi181);
not gate_53(n554,pi182);
not gate_54(n555,pi183);
not gate_55(n556,pi184);
not gate_56(n557,pi185);
not gate_57(n558,pi186);
not gate_58(n559,pi187);
not gate_59(n560,pi188);
not gate_60(n561,pi189);
not gate_61(n562,pi190);
not gate_62(n563,pi191);
not gate_63(n564,pi192);
not gate_64(n565,pi193);
not gate_65(n566,pi194);
not gate_66(n567,pi195);
not gate_67(n568,pi196);
not gate_68(n569,pi197);
not gate_69(n570,pi198);
not gate_70(n571,pi199);
not gate_71(n572,pi200);
not gate_72(n573,pi201);
not gate_73(n574,pi203);
not gate_74(n575,pi204);
not gate_75(n576,pi206);
not gate_76(n577,pi207);
not gate_77(n578,pi208);
not gate_78(n579,pi210);
not gate_79(n580,pi211);
not gate_80(n581,pi212);
not gate_81(n582,pi213);
not gate_82(n583,pi214);
not gate_83(n584,pi215);
not gate_84(n585,pi216);
not gate_85(n586,pi217);
not gate_86(n587,pi219);
not gate_87(n588,pi220);
not gate_88(n589,pi221);
not gate_89(n590,pi222);
not gate_90(n591,pi223);
not gate_91(n592,pi224);
not gate_92(n593,pi225);
not gate_93(n594,pi226);
not gate_94(n595,pi227);
not gate_95(n596,pi228);
not gate_96(n597,pi230);
not gate_97(n598,pi231);
not gate_98(n599,pi232);
not gate_99(n600,pi233);
not gate_100(n601,pi234);
not gate_101(n602,pi235);
not gate_102(n603,pi236);
not gate_103(n604,pi237);
not gate_104(n605,pi238);
not gate_105(n606,pi239);
not gate_106(n607,pi241);
not gate_107(n608,pi242);
not gate_108(n609,pi243);
not gate_109(n610,pi244);
not gate_110(n611,pi246);
not gate_111(n612,pi247);
not gate_112(n613,pi249);
not gate_113(n614,pi250);
not gate_114(n615,pi251);
not gate_115(n616,pi252);
not gate_116(n617,pi253);
not gate_117(n618,pi254);
not gate_118(n619,pi255);
and gate_119(n620,pi019,pi198);
not gate_120(n621,n620);
and gate_121(n622,pi011,n570);
not gate_122(n623,n622);
and gate_123(n624,n621,n623);
not gate_124(n625,n624);
and gate_125(n626,pi197,pi198);
not gate_126(n627,n626);
and gate_127(n628,pi195,pi196);
and gate_128(n629,n626,n628);
not gate_129(n630,n629);
and gate_130(po000,n625,n630);
and gate_131(n632,pi020,pi198);
not gate_132(n633,n632);
and gate_133(n634,pi012,n570);
not gate_134(n635,n634);
and gate_135(n636,n633,n635);
not gate_136(n637,n636);
and gate_137(po001,n630,n637);
and gate_138(n639,pi021,pi198);
not gate_139(n640,n639);
and gate_140(n641,pi013,n570);
not gate_141(n642,n641);
and gate_142(n643,n640,n642);
not gate_143(n644,n643);
and gate_144(po002,n630,n644);
and gate_145(n646,pi022,pi198);
not gate_146(n647,n646);
and gate_147(n648,pi014,n570);
not gate_148(n649,n648);
and gate_149(n650,n647,n649);
not gate_150(n651,n650);
and gate_151(po003,n630,n651);
and gate_152(n653,pi023,pi198);
not gate_153(n654,n653);
and gate_154(n655,pi015,n570);
not gate_155(n656,n655);
and gate_156(n657,n654,n656);
not gate_157(n658,n657);
and gate_158(po004,n630,n658);
and gate_159(n660,pi024,pi198);
not gate_160(n661,n660);
and gate_161(n662,pi016,n570);
not gate_162(n663,n662);
and gate_163(n664,n661,n663);
not gate_164(n665,n664);
and gate_165(po005,n630,n665);
and gate_166(n667,pi025,pi198);
not gate_167(n668,n667);
and gate_168(n669,pi017,n570);
not gate_169(n670,n669);
and gate_170(n671,n668,n670);
not gate_171(n672,n671);
and gate_172(po006,n630,n672);
and gate_173(n674,pi026,pi198);
not gate_174(n675,n674);
and gate_175(n676,pi018,n570);
not gate_176(n677,n676);
and gate_177(n678,n675,n677);
not gate_178(n679,n678);
and gate_179(po007,n630,n679);
and gate_180(n681,pi027,pi198);
not gate_181(n682,n681);
and gate_182(n683,pi019,n570);
not gate_183(n684,n683);
and gate_184(n685,n682,n684);
not gate_185(n686,n685);
and gate_186(po008,n630,n686);
and gate_187(n688,pi028,pi198);
not gate_188(n689,n688);
and gate_189(n690,pi020,n570);
not gate_190(n691,n690);
and gate_191(n692,n689,n691);
not gate_192(n693,n692);
and gate_193(po009,n630,n693);
and gate_194(n695,pi029,pi198);
not gate_195(n696,n695);
and gate_196(n697,pi021,n570);
not gate_197(n698,n697);
and gate_198(n699,n696,n698);
not gate_199(n700,n699);
and gate_200(po010,n630,n700);
and gate_201(n702,pi030,pi198);
not gate_202(n703,n702);
and gate_203(n704,pi022,n570);
not gate_204(n705,n704);
and gate_205(n706,n703,n705);
not gate_206(n707,n706);
and gate_207(po011,n630,n707);
and gate_208(n709,pi031,pi198);
not gate_209(n710,n709);
and gate_210(n711,pi023,n570);
not gate_211(n712,n711);
and gate_212(n713,n710,n712);
not gate_213(n714,n713);
and gate_214(po012,n630,n714);
and gate_215(n716,pi032,pi198);
not gate_216(n717,n716);
and gate_217(n718,pi024,n570);
not gate_218(n719,n718);
and gate_219(n720,n717,n719);
not gate_220(n721,n720);
and gate_221(po013,n630,n721);
and gate_222(n723,pi033,pi198);
not gate_223(n724,n723);
and gate_224(n725,pi025,n570);
not gate_225(n726,n725);
and gate_226(n727,n724,n726);
not gate_227(n728,n727);
and gate_228(po014,n630,n728);
and gate_229(n730,pi034,pi198);
not gate_230(n731,n730);
and gate_231(n732,pi026,n570);
not gate_232(n733,n732);
and gate_233(n734,n731,n733);
not gate_234(n735,n734);
and gate_235(po015,n630,n735);
and gate_236(n737,pi035,pi198);
not gate_237(n738,n737);
and gate_238(n739,pi027,n570);
not gate_239(n740,n739);
and gate_240(n741,n738,n740);
not gate_241(n742,n741);
and gate_242(po016,n630,n742);
and gate_243(n744,pi036,pi198);
not gate_244(n745,n744);
and gate_245(n746,pi028,n570);
not gate_246(n747,n746);
and gate_247(n748,n745,n747);
not gate_248(n749,n748);
and gate_249(po017,n630,n749);
and gate_250(n751,pi037,pi198);
not gate_251(n752,n751);
and gate_252(n753,pi029,n570);
not gate_253(n754,n753);
and gate_254(n755,n752,n754);
not gate_255(n756,n755);
and gate_256(po018,n630,n756);
and gate_257(n758,pi038,pi198);
not gate_258(n759,n758);
and gate_259(n760,pi030,n570);
not gate_260(n761,n760);
and gate_261(n762,n759,n761);
not gate_262(n763,n762);
and gate_263(po019,n630,n763);
and gate_264(n765,pi039,pi198);
not gate_265(n766,n765);
and gate_266(n767,pi031,n570);
not gate_267(n768,n767);
and gate_268(n769,n766,n768);
not gate_269(n770,n769);
and gate_270(po020,n630,n770);
and gate_271(n772,pi040,pi198);
not gate_272(n773,n772);
and gate_273(n774,pi032,n570);
not gate_274(n775,n774);
and gate_275(n776,n773,n775);
not gate_276(n777,n776);
and gate_277(po021,n630,n777);
and gate_278(n779,pi041,pi198);
not gate_279(n780,n779);
and gate_280(n781,pi033,n570);
not gate_281(n782,n781);
and gate_282(n783,n780,n782);
not gate_283(n784,n783);
and gate_284(po022,n630,n784);
and gate_285(n786,pi042,pi198);
not gate_286(n787,n786);
and gate_287(n788,pi034,n570);
not gate_288(n789,n788);
and gate_289(n790,n787,n789);
not gate_290(n791,n790);
and gate_291(po023,n630,n791);
and gate_292(n793,pi043,pi198);
not gate_293(n794,n793);
and gate_294(n795,pi035,n570);
not gate_295(n796,n795);
and gate_296(n797,n794,n796);
not gate_297(n798,n797);
and gate_298(po024,n630,n798);
and gate_299(n800,pi044,pi198);
not gate_300(n801,n800);
and gate_301(n802,pi036,n570);
not gate_302(n803,n802);
and gate_303(n804,n801,n803);
not gate_304(n805,n804);
and gate_305(po025,n630,n805);
and gate_306(n807,pi045,pi198);
not gate_307(n808,n807);
and gate_308(n809,pi037,n570);
not gate_309(n810,n809);
and gate_310(n811,n808,n810);
not gate_311(n812,n811);
and gate_312(po026,n630,n812);
and gate_313(n814,pi046,pi198);
not gate_314(n815,n814);
and gate_315(n816,pi038,n570);
not gate_316(n817,n816);
and gate_317(n818,n815,n817);
not gate_318(n819,n818);
and gate_319(po027,n630,n819);
and gate_320(n821,pi047,pi198);
not gate_321(n822,n821);
and gate_322(n823,pi039,n570);
not gate_323(n824,n823);
and gate_324(n825,n822,n824);
not gate_325(n826,n825);
and gate_326(po028,n630,n826);
and gate_327(n828,pi048,pi198);
not gate_328(n829,n828);
and gate_329(n830,pi040,n570);
not gate_330(n831,n830);
and gate_331(n832,n829,n831);
not gate_332(n833,n832);
and gate_333(po029,n630,n833);
and gate_334(n835,pi049,pi198);
not gate_335(n836,n835);
and gate_336(n837,pi041,n570);
not gate_337(n838,n837);
and gate_338(n839,n836,n838);
not gate_339(n840,n839);
and gate_340(po030,n630,n840);
and gate_341(n842,pi050,pi198);
not gate_342(n843,n842);
and gate_343(n844,pi042,n570);
not gate_344(n845,n844);
and gate_345(n846,n843,n845);
not gate_346(n847,n846);
and gate_347(po031,n630,n847);
and gate_348(n849,pi051,pi198);
not gate_349(n850,n849);
and gate_350(n851,pi043,n570);
not gate_351(n852,n851);
and gate_352(n853,n850,n852);
not gate_353(n854,n853);
and gate_354(po032,n630,n854);
and gate_355(n856,pi052,pi198);
not gate_356(n857,n856);
and gate_357(n858,pi044,n570);
not gate_358(n859,n858);
and gate_359(n860,n857,n859);
not gate_360(n861,n860);
and gate_361(po033,n630,n861);
and gate_362(n863,pi053,pi198);
not gate_363(n864,n863);
and gate_364(n865,pi045,n570);
not gate_365(n866,n865);
and gate_366(n867,n864,n866);
not gate_367(n868,n867);
and gate_368(po034,n630,n868);
and gate_369(n870,pi054,pi198);
not gate_370(n871,n870);
and gate_371(n872,pi046,n570);
not gate_372(n873,n872);
and gate_373(n874,n871,n873);
not gate_374(n875,n874);
and gate_375(po035,n630,n875);
and gate_376(n877,pi055,pi198);
not gate_377(n878,n877);
and gate_378(n879,pi047,n570);
not gate_379(n880,n879);
and gate_380(n881,n878,n880);
not gate_381(n882,n881);
and gate_382(po036,n630,n882);
and gate_383(n884,pi056,pi198);
not gate_384(n885,n884);
and gate_385(n886,pi048,n570);
not gate_386(n887,n886);
and gate_387(n888,n885,n887);
not gate_388(n889,n888);
and gate_389(po037,n630,n889);
and gate_390(n891,pi049,n570);
not gate_391(n892,n891);
and gate_392(n893,pi057,pi198);
not gate_393(n894,n893);
and gate_394(n895,n892,n894);
not gate_395(n896,n895);
and gate_396(po038,n630,n896);
and gate_397(n898,pi050,n570);
not gate_398(n899,n898);
and gate_399(n900,pi058,pi198);
not gate_400(n901,n900);
and gate_401(n902,n899,n901);
not gate_402(n903,n902);
and gate_403(po039,n630,n903);
and gate_404(n905,pi051,n570);
not gate_405(n906,n905);
and gate_406(n907,pi059,pi198);
not gate_407(n908,n907);
and gate_408(n909,n906,n908);
not gate_409(n910,n909);
and gate_410(po040,n630,n910);
and gate_411(n912,pi052,n570);
not gate_412(n913,n912);
and gate_413(n914,pi060,pi198);
not gate_414(n915,n914);
and gate_415(n916,n913,n915);
not gate_416(n917,n916);
and gate_417(po041,n630,n917);
and gate_418(n919,pi053,n570);
not gate_419(n920,n919);
and gate_420(n921,pi061,pi198);
not gate_421(n922,n921);
and gate_422(n923,n920,n922);
not gate_423(n924,n923);
and gate_424(po042,n630,n924);
and gate_425(n926,pi054,n570);
not gate_426(n927,n926);
and gate_427(n928,pi062,pi198);
not gate_428(n929,n928);
and gate_429(n930,n927,n929);
not gate_430(n931,n930);
and gate_431(po043,n630,n931);
and gate_432(n933,pi055,n570);
not gate_433(n934,n933);
and gate_434(n935,pi063,pi198);
not gate_435(n936,n935);
and gate_436(n937,n934,n936);
not gate_437(n938,n937);
and gate_438(po044,n630,n938);
and gate_439(n940,pi056,n570);
not gate_440(n941,n940);
and gate_441(n942,pi064,pi198);
not gate_442(n943,n942);
and gate_443(n944,n941,n943);
not gate_444(n945,n944);
and gate_445(po045,n630,n945);
and gate_446(n947,pi065,pi198);
not gate_447(n948,n947);
and gate_448(n949,pi057,n570);
not gate_449(n950,n949);
and gate_450(n951,n948,n950);
not gate_451(n952,n951);
and gate_452(po046,n630,n952);
and gate_453(n954,pi066,pi198);
not gate_454(n955,n954);
and gate_455(n956,pi058,n570);
not gate_456(n957,n956);
and gate_457(n958,n955,n957);
not gate_458(n959,n958);
and gate_459(po047,n630,n959);
and gate_460(n961,pi000,pi198);
not gate_461(n962,n961);
and gate_462(n963,pi059,n570);
not gate_463(n964,n963);
and gate_464(n965,n962,n964);
not gate_465(n966,n965);
and gate_466(po048,n630,n966);
and gate_467(n968,pi001,pi198);
not gate_468(n969,n968);
and gate_469(n970,pi060,n570);
not gate_470(n971,n970);
and gate_471(n972,n969,n971);
not gate_472(n973,n972);
and gate_473(po049,n630,n973);
and gate_474(n975,pi002,pi198);
not gate_475(n976,n975);
and gate_476(n977,pi061,n570);
not gate_477(n978,n977);
and gate_478(n979,n976,n978);
not gate_479(n980,n979);
and gate_480(po050,n630,n980);
and gate_481(n982,pi003,pi198);
not gate_482(n983,n982);
and gate_483(n984,pi062,n570);
not gate_484(n985,n984);
and gate_485(n986,n983,n985);
not gate_486(n987,n986);
and gate_487(po051,n630,n987);
and gate_488(n989,pi004,pi198);
not gate_489(n990,n989);
and gate_490(n991,pi063,n570);
not gate_491(n992,n991);
and gate_492(n993,n990,n992);
not gate_493(n994,n993);
and gate_494(po052,n630,n994);
and gate_495(n996,pi005,pi198);
not gate_496(n997,n996);
and gate_497(n998,pi064,n570);
not gate_498(n999,n998);
and gate_499(n1000,n997,n999);
not gate_500(n1001,n1000);
and gate_501(po053,n630,n1001);
and gate_502(n1003,pi006,pi198);
not gate_503(n1004,n1003);
and gate_504(n1005,pi065,n570);
not gate_505(n1006,n1005);
and gate_506(n1007,n1004,n1006);
not gate_507(n1008,n1007);
and gate_508(po054,n630,n1008);
and gate_509(n1010,pi007,pi198);
not gate_510(n1011,n1010);
and gate_511(n1012,pi066,n570);
not gate_512(n1013,n1012);
and gate_513(n1014,n1011,n1013);
not gate_514(n1015,n1014);
and gate_515(po055,n630,n1015);
and gate_516(n1017,pi142,n596);
not gate_517(n1018,n1017);
and gate_518(n1019,n514,pi228);
not gate_519(n1020,n1019);
and gate_520(n1021,n1018,n1020);
not gate_521(n1022,n1021);
and gate_522(n1023,pi143,n603);
not gate_523(n1024,n1023);
and gate_524(n1025,n515,pi236);
not gate_525(n1026,n1025);
and gate_526(n1027,n1024,n1026);
not gate_527(n1028,n1027);
and gate_528(n1029,pi144,n611);
not gate_529(n1030,n1029);
and gate_530(n1031,n516,pi246);
not gate_531(n1032,n1031);
and gate_532(n1033,n1030,n1032);
not gate_533(n1034,n1033);
and gate_534(n1035,pi145,n616);
not gate_535(n1036,n1035);
and gate_536(n1037,n517,pi252);
not gate_537(n1038,n1037);
and gate_538(n1039,n1036,n1038);
not gate_539(n1040,n1039);
and gate_540(n1041,pi147,n608);
not gate_541(n1042,n1041);
and gate_542(n1043,n519,pi242);
not gate_543(n1044,n1043);
and gate_544(n1045,n1042,n1044);
not gate_545(n1046,n1045);
and gate_546(n1047,pi146,n598);
not gate_547(n1048,n1047);
and gate_548(n1049,n518,pi231);
not gate_549(n1050,n1049);
and gate_550(n1051,n1048,n1050);
not gate_551(n1052,n1051);
and gate_552(n1053,n1045,n1051);
and gate_553(n1054,n1040,n1053);
and gate_554(n1055,n1033,n1054);
and gate_555(n1056,n1028,n1055);
and gate_556(n1057,n1021,n1056);
not gate_557(n1058,n1057);
and gate_558(n1059,n1034,n1054);
and gate_559(n1060,n1027,n1059);
and gate_560(n1061,n1021,n1060);
not gate_561(n1062,n1061);
and gate_562(n1063,n1058,n1062);
and gate_563(n1064,n1021,n1027);
and gate_564(n1065,n1055,n1064);
not gate_565(n1066,n1065);
and gate_566(n1067,n1063,n1066);
and gate_567(n1068,n1021,n1028);
and gate_568(n1069,n1059,n1068);
not gate_569(n1070,n1069);
and gate_570(n1071,n1045,n1052);
and gate_571(n1072,n1040,n1071);
and gate_572(n1073,n1034,n1072);
and gate_573(n1074,n1064,n1073);
not gate_574(n1075,n1074);
and gate_575(n1076,n1070,n1075);
and gate_576(n1077,n1039,n1071);
and gate_577(n1078,n1034,n1077);
and gate_578(n1079,n1021,n1078);
not gate_579(n1080,n1079);
and gate_580(n1081,n1076,n1080);
and gate_581(n1082,n1067,n1081);
and gate_582(n1083,n1039,n1051);
and gate_583(n1084,n1045,n1083);
and gate_584(n1085,n1033,n1084);
and gate_585(n1086,n1028,n1085);
and gate_586(n1087,n1022,n1086);
not gate_587(n1088,n1087);
and gate_588(n1089,n1022,n1056);
not gate_589(n1090,n1089);
and gate_590(n1091,n1088,n1090);
and gate_591(n1092,n1022,n1027);
and gate_592(n1093,n1085,n1092);
not gate_593(n1094,n1093);
and gate_594(n1095,n1091,n1094);
and gate_595(n1096,n1027,n1078);
and gate_596(n1097,n1022,n1096);
not gate_597(n1098,n1097);
and gate_598(n1099,n1028,n1073);
and gate_599(n1100,n1022,n1099);
not gate_600(n1101,n1100);
and gate_601(n1102,n1098,n1101);
and gate_602(n1103,n1028,n1078);
and gate_603(n1104,n1022,n1103);
not gate_604(n1105,n1104);
and gate_605(n1106,n1033,n1072);
and gate_606(n1107,n1027,n1106);
and gate_607(n1108,n1022,n1107);
not gate_608(n1109,n1108);
and gate_609(n1110,n1105,n1109);
and gate_610(n1111,n1102,n1110);
and gate_611(n1112,n1095,n1111);
and gate_612(n1113,n1082,n1112);
and gate_613(n1114,n1046,n1051);
and gate_614(n1115,n1039,n1114);
and gate_615(n1116,n1034,n1115);
and gate_616(n1117,n1028,n1116);
and gate_617(n1118,n1021,n1117);
not gate_618(n1119,n1118);
and gate_619(n1120,n1040,n1114);
and gate_620(n1121,n1033,n1120);
and gate_621(n1122,n1064,n1121);
not gate_622(n1123,n1122);
and gate_623(n1124,n1034,n1120);
and gate_624(n1125,n1064,n1124);
not gate_625(n1126,n1125);
and gate_626(n1127,n1123,n1126);
and gate_627(n1128,n1119,n1127);
and gate_628(n1129,n1046,n1052);
and gate_629(n1130,n1040,n1129);
and gate_630(n1131,n1033,n1130);
and gate_631(n1132,n1027,n1131);
and gate_632(n1133,n1021,n1132);
not gate_633(n1134,n1133);
and gate_634(n1135,n1034,n1130);
and gate_635(n1136,n1028,n1135);
and gate_636(n1137,n1021,n1136);
not gate_637(n1138,n1137);
and gate_638(n1139,n1134,n1138);
and gate_639(n1140,n1039,n1129);
and gate_640(n1141,n1033,n1140);
and gate_641(n1142,n1027,n1141);
and gate_642(n1143,n1021,n1142);
not gate_643(n1144,n1143);
and gate_644(n1145,n1068,n1131);
not gate_645(n1146,n1145);
and gate_646(n1147,n1144,n1146);
and gate_647(n1148,n1139,n1147);
and gate_648(n1149,n1128,n1148);
and gate_649(n1150,n1022,n1117);
not gate_650(n1151,n1150);
and gate_651(n1152,n1028,n1121);
and gate_652(n1153,n1022,n1152);
not gate_653(n1154,n1153);
and gate_654(n1155,n1151,n1154);
and gate_655(n1156,n1022,n1033);
and gate_656(n1157,n1027,n1115);
and gate_657(n1158,n1156,n1157);
not gate_658(n1159,n1158);
and gate_659(n1160,n1155,n1159);
and gate_660(n1161,n1022,n1132);
not gate_661(n1162,n1161);
and gate_662(n1163,n1022,n1136);
not gate_663(n1164,n1163);
and gate_664(n1165,n1162,n1164);
and gate_665(n1166,n1022,n1141);
not gate_666(n1167,n1166);
and gate_667(n1168,n1165,n1167);
and gate_668(n1169,n1160,n1168);
and gate_669(n1170,n1149,n1169);
and gate_670(n1171,n1113,n1170);
and gate_671(n1172,n1040,n1092);
and gate_672(n1173,n1034,n1172);
not gate_673(n1174,n1173);
and gate_674(n1175,n1021,n1033);
not gate_675(n1176,n1175);
and gate_676(n1177,n1039,n1175);
and gate_677(n1178,n1028,n1177);
not gate_678(n1179,n1178);
and gate_679(n1180,n1174,n1179);
not gate_680(n1181,n1180);
and gate_681(n1182,n1046,n1181);
not gate_682(n1183,n1182);
and gate_683(n1184,n1022,n1034);
not gate_684(n1185,n1184);
and gate_685(n1186,n1176,n1185);
not gate_686(n1187,n1186);
and gate_687(n1188,n1027,n1187);
and gate_688(n1189,n1039,n1188);
and gate_689(n1190,n1045,n1189);
not gate_690(n1191,n1190);
and gate_691(n1192,n1183,n1191);
not gate_692(n1193,n1192);
and gate_693(n1194,n1051,n1193);
not gate_694(n1195,n1194);
and gate_695(n1196,n1171,n1195);
not gate_696(n1197,n1196);
and gate_697(n1198,n542,n1197);
not gate_698(n1199,n1198);
and gate_699(n1200,pi170,n1196);
not gate_700(n1201,n1200);
and gate_701(n1202,n1199,n1201);
not gate_702(n1203,n1202);
and gate_703(n1204,n629,n1203);
not gate_704(n1205,n1204);
and gate_705(n1206,pi067,n570);
not gate_706(n1207,n1206);
and gate_707(n1208,n1205,n1207);
not gate_708(po056,n1208);
and gate_709(n1210,pi138,n629);
not gate_710(n1211,n1210);
and gate_711(n1212,pi068,n570);
not gate_712(n1213,n1212);
and gate_713(n1214,n1211,n1213);
not gate_714(po057,n1214);
and gate_715(n1216,pi158,n590);
not gate_716(n1217,n1216);
and gate_717(n1218,n530,pi222);
not gate_718(n1219,n1218);
and gate_719(n1220,n1217,n1219);
not gate_720(n1221,n1220);
and gate_721(n1222,pi159,n594);
not gate_722(n1223,n1222);
and gate_723(n1224,n531,pi226);
not gate_724(n1225,n1224);
and gate_725(n1226,n1223,n1225);
not gate_726(n1227,n1226);
and gate_727(n1228,pi160,n574);
not gate_728(n1229,n1228);
and gate_729(n1230,n532,pi203);
not gate_730(n1231,n1230);
and gate_731(n1232,n1229,n1231);
not gate_732(n1233,n1232);
and gate_733(n1234,pi161,n585);
not gate_734(n1235,n1234);
and gate_735(n1236,n533,pi216);
not gate_736(n1237,n1236);
and gate_737(n1238,n1235,n1237);
not gate_738(n1239,n1238);
and gate_739(n1240,pi131,n582);
not gate_740(n1241,n1240);
and gate_741(n1242,n503,pi213);
not gate_742(n1243,n1242);
and gate_743(n1244,n1241,n1243);
not gate_744(n1245,n1244);
and gate_745(n1246,pi162,n579);
not gate_746(n1247,n1246);
and gate_747(n1248,n534,pi210);
not gate_748(n1249,n1248);
and gate_749(n1250,n1247,n1249);
not gate_750(n1251,n1250);
and gate_751(n1252,n1244,n1251);
and gate_752(n1253,n1238,n1252);
and gate_753(n1254,n1233,n1253);
and gate_754(n1255,n1226,n1254);
and gate_755(n1256,n1220,n1255);
not gate_756(n1257,n1256);
and gate_757(n1258,n1227,n1254);
and gate_758(n1259,n1220,n1258);
not gate_759(n1260,n1259);
and gate_760(n1261,n1257,n1260);
and gate_761(n1262,n1244,n1250);
and gate_762(n1263,n1238,n1262);
and gate_763(n1264,n1232,n1263);
and gate_764(n1265,n1220,n1226);
not gate_765(n1266,n1265);
and gate_766(n1267,n1264,n1265);
not gate_767(n1268,n1267);
and gate_768(n1269,n1261,n1268);
and gate_769(n1270,n1239,n1252);
and gate_770(n1271,n1232,n1270);
and gate_771(n1272,n1226,n1271);
and gate_772(n1273,n1220,n1272);
not gate_773(n1274,n1273);
and gate_774(n1275,n1233,n1270);
and gate_775(n1276,n1220,n1227);
and gate_776(n1277,n1275,n1276);
not gate_777(n1278,n1277);
and gate_778(n1279,n1274,n1278);
and gate_779(n1280,n1233,n1263);
and gate_780(n1281,n1226,n1280);
and gate_781(n1282,n1221,n1281);
not gate_782(n1283,n1282);
and gate_783(n1284,n1221,n1227);
not gate_784(n1285,n1284);
and gate_785(n1286,n1264,n1284);
not gate_786(n1287,n1286);
and gate_787(n1288,n1283,n1287);
and gate_788(n1289,n1279,n1288);
and gate_789(n1290,n1269,n1289);
and gate_790(n1291,n1239,n1262);
and gate_791(n1292,n1233,n1291);
and gate_792(n1293,n1226,n1292);
and gate_793(n1294,n1221,n1293);
not gate_794(n1295,n1294);
and gate_795(n1296,n1232,n1253);
and gate_796(n1297,n1227,n1296);
and gate_797(n1298,n1221,n1297);
not gate_798(n1299,n1298);
and gate_799(n1300,n1295,n1299);
and gate_800(n1301,n1232,n1291);
and gate_801(n1302,n1221,n1226);
and gate_802(n1303,n1301,n1302);
not gate_803(n1304,n1303);
and gate_804(n1305,n1300,n1304);
and gate_805(n1306,n1221,n1255);
not gate_806(n1307,n1306);
and gate_807(n1308,n1227,n1271);
and gate_808(n1309,n1221,n1308);
not gate_809(n1310,n1309);
and gate_810(n1311,n1307,n1310);
and gate_811(n1312,n1220,n1281);
not gate_812(n1313,n1312);
and gate_813(n1314,n1245,n1250);
and gate_814(n1315,n1238,n1314);
and gate_815(n1316,n1233,n1315);
and gate_816(n1317,n1265,n1316);
not gate_817(n1318,n1317);
and gate_818(n1319,n1313,n1318);
and gate_819(n1320,n1311,n1319);
and gate_820(n1321,n1305,n1320);
and gate_821(n1322,n1290,n1321);
and gate_822(n1323,n1239,n1314);
and gate_823(n1324,n1232,n1323);
and gate_824(n1325,n1227,n1324);
and gate_825(n1326,n1220,n1325);
not gate_826(n1327,n1326);
and gate_827(n1328,n1245,n1251);
and gate_828(n1329,n1238,n1328);
and gate_829(n1330,n1232,n1329);
and gate_830(n1331,n1226,n1330);
and gate_831(n1332,n1220,n1331);
not gate_832(n1333,n1332);
and gate_833(n1334,n1327,n1333);
and gate_834(n1335,n1265,n1324);
not gate_835(n1336,n1335);
and gate_836(n1337,n1334,n1336);
and gate_837(n1338,n1227,n1330);
and gate_838(n1339,n1220,n1338);
not gate_839(n1340,n1339);
and gate_840(n1341,n1233,n1329);
and gate_841(n1342,n1227,n1341);
and gate_842(n1343,n1220,n1342);
not gate_843(n1344,n1343);
and gate_844(n1345,n1340,n1344);
and gate_845(n1346,n1239,n1328);
and gate_846(n1347,n1233,n1346);
and gate_847(n1348,n1226,n1347);
and gate_848(n1349,n1220,n1348);
not gate_849(n1350,n1349);
and gate_850(n1351,n1232,n1315);
and gate_851(n1352,n1302,n1351);
not gate_852(n1353,n1352);
and gate_853(n1354,n1350,n1353);
and gate_854(n1355,n1345,n1354);
and gate_855(n1356,n1337,n1355);
and gate_856(n1357,n1233,n1323);
and gate_857(n1358,n1227,n1357);
and gate_858(n1359,n1221,n1358);
not gate_859(n1360,n1359);
and gate_860(n1361,n1221,n1331);
not gate_861(n1362,n1361);
and gate_862(n1363,n1360,n1362);
and gate_863(n1364,n1284,n1351);
not gate_864(n1365,n1364);
and gate_865(n1366,n1363,n1365);
and gate_866(n1367,n1221,n1342);
not gate_867(n1368,n1367);
and gate_868(n1369,n1276,n1301);
not gate_869(n1370,n1369);
and gate_870(n1371,n1368,n1370);
and gate_871(n1372,n1221,n1348);
not gate_872(n1373,n1372);
and gate_873(n1374,n1284,n1347);
not gate_874(n1375,n1374);
and gate_875(n1376,n1373,n1375);
and gate_876(n1377,n1371,n1376);
and gate_877(n1378,n1366,n1377);
and gate_878(n1379,n1356,n1378);
and gate_879(n1380,n1322,n1379);
and gate_880(n1381,n1221,n1239);
not gate_881(n1382,n1381);
and gate_882(n1383,n1220,n1238);
not gate_883(n1384,n1383);
and gate_884(n1385,n1382,n1384);
not gate_885(n1386,n1385);
and gate_886(n1387,n1226,n1386);
and gate_887(n1388,n1245,n1387);
not gate_888(n1389,n1388);
and gate_889(n1390,n1238,n1244);
not gate_890(n1391,n1390);
and gate_891(n1392,n1276,n1390);
not gate_892(n1393,n1392);
and gate_893(n1394,n1389,n1393);
not gate_894(n1395,n1394);
and gate_895(n1396,n1232,n1395);
not gate_896(n1397,n1396);
and gate_897(n1398,n1233,n1284);
and gate_898(n1399,n1390,n1398);
not gate_899(n1400,n1399);
and gate_900(n1401,n1397,n1400);
not gate_901(n1402,n1401);
and gate_902(n1403,n1250,n1402);
not gate_903(n1404,n1403);
and gate_904(n1405,n1380,n1404);
not gate_905(n1406,n1405);
and gate_906(n1407,n550,n1406);
not gate_907(n1408,n1407);
and gate_908(n1409,pi178,n1405);
not gate_909(n1410,n1409);
and gate_910(n1411,n1408,n1410);
not gate_911(n1412,n1411);
and gate_912(n1413,n629,n1412);
not gate_913(n1414,n1413);
and gate_914(n1415,pi069,n570);
not gate_915(n1416,n1415);
and gate_916(n1417,n1414,n1416);
not gate_917(po058,n1417);
and gate_918(n1419,pi146,n629);
not gate_919(n1420,n1419);
and gate_920(n1421,pi070,n570);
not gate_921(n1422,n1421);
and gate_922(n1423,n1420,n1422);
not gate_923(po059,n1423);
and gate_924(n1425,n1220,n1308);
not gate_925(n1426,n1425);
and gate_926(n1427,n1260,n1426);
and gate_927(n1428,n1268,n1427);
and gate_928(n1429,n1226,n1296);
and gate_929(n1430,n1221,n1429);
not gate_930(n1431,n1430);
and gate_931(n1432,n1304,n1431);
and gate_932(n1433,n1287,n1295);
and gate_933(n1434,n1432,n1433);
and gate_934(n1435,n1428,n1434);
and gate_935(n1436,n1221,n1258);
not gate_936(n1437,n1436);
and gate_937(n1438,n1221,n1272);
not gate_938(n1439,n1438);
and gate_939(n1440,n1437,n1439);
and gate_940(n1441,n1307,n1440);
and gate_941(n1442,n1220,n1358);
not gate_942(n1443,n1442);
and gate_943(n1444,n1336,n1443);
and gate_944(n1445,n1319,n1444);
and gate_945(n1446,n1441,n1445);
and gate_946(n1447,n1435,n1446);
and gate_947(n1448,n1226,n1341);
and gate_948(n1449,n1220,n1448);
not gate_949(n1450,n1449);
and gate_950(n1451,n1340,n1450);
and gate_951(n1452,n1333,n1451);
and gate_952(n1453,n1232,n1346);
and gate_953(n1454,n1276,n1453);
not gate_954(n1455,n1454);
and gate_955(n1456,n1353,n1455);
and gate_956(n1457,n1221,n1325);
not gate_957(n1458,n1457);
and gate_958(n1459,n1365,n1458);
and gate_959(n1460,n1456,n1459);
and gate_960(n1461,n1452,n1460);
and gate_961(n1462,n1221,n1338);
not gate_962(n1463,n1462);
and gate_963(n1464,n1371,n1463);
and gate_964(n1465,n1226,n1453);
and gate_965(n1466,n1221,n1465);
not gate_966(n1467,n1466);
and gate_967(n1468,n1375,n1467);
and gate_968(n1469,n1220,n1293);
not gate_969(n1470,n1469);
and gate_970(n1471,n1220,n1297);
not gate_971(n1472,n1471);
and gate_972(n1473,n1470,n1472);
and gate_973(n1474,n1468,n1473);
and gate_974(n1475,n1464,n1474);
and gate_975(n1476,n1461,n1475);
and gate_976(n1477,n1447,n1476);
and gate_977(n1478,n1266,n1285);
not gate_978(n1479,n1478);
and gate_979(n1480,n1238,n1478);
not gate_980(n1481,n1480);
and gate_981(n1482,n1244,n1276);
not gate_982(n1483,n1482);
and gate_983(n1484,n1481,n1483);
not gate_984(n1485,n1484);
and gate_985(n1486,n1391,n1485);
and gate_986(n1487,n1250,n1486);
not gate_987(n1488,n1487);
and gate_988(n1489,n1270,n1284);
not gate_989(n1490,n1489);
and gate_990(n1491,n1488,n1490);
not gate_991(n1492,n1491);
and gate_992(n1493,n1233,n1492);
not gate_993(n1494,n1493);
and gate_994(n1495,n1477,n1494);
not gate_995(n1496,n1495);
and gate_996(n1497,n558,n1496);
not gate_997(n1498,n1497);
and gate_998(n1499,pi186,n1495);
not gate_999(n1500,n1499);
and gate_1000(n1501,n1498,n1500);
not gate_1001(n1502,n1501);
and gate_1002(n1503,n629,n1502);
not gate_1003(n1504,n1503);
and gate_1004(n1505,pi071,n570);
not gate_1005(n1506,n1505);
and gate_1006(n1507,n1504,n1506);
not gate_1007(po060,n1507);
and gate_1008(n1509,pi154,n629);
not gate_1009(n1510,n1509);
and gate_1010(n1511,pi072,n570);
not gate_1011(n1512,n1511);
and gate_1012(n1513,n1510,n1512);
not gate_1013(po061,n1513);
and gate_1014(n1515,pi146,n593);
not gate_1015(n1516,n1515);
and gate_1016(n1517,n518,pi225);
not gate_1017(n1518,n1517);
and gate_1018(n1519,n1516,n1518);
not gate_1019(n1520,n1519);
and gate_1020(n1521,pi147,n583);
not gate_1021(n1522,n1521);
and gate_1022(n1523,n519,pi214);
not gate_1023(n1524,n1523);
and gate_1024(n1525,n1522,n1524);
not gate_1025(n1526,n1525);
and gate_1026(n1527,pi148,n577);
not gate_1027(n1528,n1527);
and gate_1028(n1529,n520,pi207);
not gate_1029(n1530,n1529);
and gate_1030(n1531,n1528,n1530);
not gate_1031(n1532,n1531);
and gate_1032(n1533,pi149,n572);
not gate_1033(n1534,n1533);
and gate_1034(n1535,n521,pi200);
not gate_1035(n1536,n1535);
and gate_1036(n1537,n1534,n1536);
not gate_1037(n1538,n1537);
and gate_1038(n1539,pi151,n580);
not gate_1039(n1540,n1539);
and gate_1040(n1541,n523,pi211);
not gate_1041(n1542,n1541);
and gate_1042(n1543,n1540,n1542);
not gate_1043(n1544,n1543);
and gate_1044(n1545,pi150,n588);
not gate_1045(n1546,n1545);
and gate_1046(n1547,n522,pi220);
not gate_1047(n1548,n1547);
and gate_1048(n1549,n1546,n1548);
not gate_1049(n1550,n1549);
and gate_1050(n1551,n1543,n1549);
and gate_1051(n1552,n1537,n1551);
and gate_1052(n1553,n1531,n1552);
and gate_1053(n1554,n1525,n1553);
and gate_1054(n1555,n1519,n1554);
not gate_1055(n1556,n1555);
and gate_1056(n1557,n1532,n1552);
and gate_1057(n1558,n1526,n1557);
and gate_1058(n1559,n1519,n1558);
not gate_1059(n1560,n1559);
and gate_1060(n1561,n1519,n1526);
and gate_1061(n1562,n1553,n1561);
not gate_1062(n1563,n1562);
and gate_1063(n1564,n1560,n1563);
and gate_1064(n1565,n1556,n1564);
and gate_1065(n1566,n1543,n1550);
and gate_1066(n1567,n1537,n1566);
and gate_1067(n1568,n1532,n1567);
and gate_1068(n1569,n1526,n1568);
and gate_1069(n1570,n1519,n1569);
not gate_1070(n1571,n1570);
and gate_1071(n1572,n1538,n1551);
and gate_1072(n1573,n1532,n1572);
and gate_1073(n1574,n1519,n1525);
and gate_1074(n1575,n1573,n1574);
not gate_1075(n1576,n1575);
and gate_1076(n1577,n1571,n1576);
and gate_1077(n1578,n1538,n1566);
and gate_1078(n1579,n1532,n1578);
and gate_1079(n1580,n1526,n1579);
and gate_1080(n1581,n1519,n1580);
not gate_1081(n1582,n1581);
and gate_1082(n1583,n1531,n1578);
and gate_1083(n1584,n1574,n1583);
not gate_1084(n1585,n1584);
and gate_1085(n1586,n1582,n1585);
and gate_1086(n1587,n1577,n1586);
and gate_1087(n1588,n1565,n1587);
and gate_1088(n1589,n1520,n1554);
not gate_1089(n1590,n1589);
and gate_1090(n1591,n1525,n1557);
and gate_1091(n1592,n1520,n1591);
not gate_1092(n1593,n1592);
and gate_1093(n1594,n1520,n1558);
not gate_1094(n1595,n1594);
and gate_1095(n1596,n1593,n1595);
and gate_1096(n1597,n1590,n1596);
and gate_1097(n1598,n1531,n1572);
and gate_1098(n1599,n1526,n1598);
and gate_1099(n1600,n1520,n1599);
not gate_1100(n1601,n1600);
and gate_1101(n1602,n1520,n1526);
and gate_1102(n1603,n1531,n1602);
and gate_1103(n1604,n1567,n1603);
not gate_1104(n1605,n1604);
and gate_1105(n1606,n1601,n1605);
and gate_1106(n1607,n1526,n1573);
and gate_1107(n1608,n1520,n1607);
not gate_1108(n1609,n1608);
and gate_1109(n1610,n1520,n1580);
not gate_1110(n1611,n1610);
and gate_1111(n1612,n1609,n1611);
and gate_1112(n1613,n1606,n1612);
and gate_1113(n1614,n1597,n1613);
and gate_1114(n1615,n1588,n1614);
and gate_1115(n1616,n1544,n1549);
and gate_1116(n1617,n1538,n1616);
and gate_1117(n1618,n1532,n1617);
and gate_1118(n1619,n1525,n1618);
and gate_1119(n1620,n1519,n1619);
not gate_1120(n1621,n1620);
and gate_1121(n1622,n1531,n1617);
and gate_1122(n1623,n1561,n1622);
not gate_1123(n1624,n1623);
and gate_1124(n1625,n1621,n1624);
and gate_1125(n1626,n1537,n1616);
and gate_1126(n1627,n1532,n1626);
and gate_1127(n1628,n1574,n1627);
not gate_1128(n1629,n1628);
and gate_1129(n1630,n1625,n1629);
and gate_1130(n1631,n1544,n1550);
and gate_1131(n1632,n1537,n1631);
and gate_1132(n1633,n1531,n1632);
and gate_1133(n1634,n1525,n1633);
and gate_1134(n1635,n1519,n1634);
not gate_1135(n1636,n1635);
and gate_1136(n1637,n1561,n1618);
not gate_1137(n1638,n1637);
and gate_1138(n1639,n1636,n1638);
and gate_1139(n1640,n1532,n1632);
and gate_1140(n1641,n1525,n1640);
and gate_1141(n1642,n1519,n1641);
not gate_1142(n1643,n1642);
and gate_1143(n1644,n1538,n1631);
and gate_1144(n1645,n1531,n1644);
and gate_1145(n1646,n1525,n1645);
and gate_1146(n1647,n1519,n1646);
not gate_1147(n1648,n1647);
and gate_1148(n1649,n1643,n1648);
and gate_1149(n1650,n1639,n1649);
and gate_1150(n1651,n1630,n1650);
and gate_1151(n1652,n1531,n1626);
and gate_1152(n1653,n1525,n1652);
and gate_1153(n1654,n1520,n1653);
not gate_1154(n1655,n1654);
and gate_1155(n1656,n1526,n1652);
and gate_1156(n1657,n1520,n1656);
not gate_1157(n1658,n1657);
and gate_1158(n1659,n1520,n1619);
not gate_1159(n1660,n1659);
and gate_1160(n1661,n1658,n1660);
and gate_1161(n1662,n1655,n1661);
and gate_1162(n1663,n1520,n1634);
not gate_1163(n1664,n1663);
and gate_1164(n1665,n1520,n1641);
not gate_1165(n1666,n1665);
and gate_1166(n1667,n1664,n1666);
and gate_1167(n1668,n1526,n1640);
and gate_1168(n1669,n1520,n1668);
not gate_1169(n1670,n1669);
and gate_1170(n1671,n1602,n1645);
not gate_1171(n1672,n1671);
and gate_1172(n1673,n1670,n1672);
and gate_1173(n1674,n1667,n1673);
and gate_1174(n1675,n1662,n1674);
and gate_1175(n1676,n1651,n1675);
and gate_1176(n1677,n1615,n1676);
and gate_1177(n1678,n1520,n1538);
not gate_1178(n1679,n1678);
and gate_1179(n1680,n1549,n1678);
not gate_1180(n1681,n1680);
and gate_1181(n1682,n1519,n1537);
not gate_1182(n1683,n1682);
and gate_1183(n1684,n1550,n1682);
not gate_1184(n1685,n1684);
and gate_1185(n1686,n1681,n1685);
not gate_1186(n1687,n1686);
and gate_1187(n1688,n1526,n1544);
not gate_1188(n1689,n1688);
and gate_1189(n1690,n1687,n1688);
not gate_1190(n1691,n1690);
and gate_1191(n1692,n1679,n1683);
not gate_1192(n1693,n1692);
and gate_1193(n1694,n1525,n1693);
and gate_1194(n1695,n1566,n1694);
not gate_1195(n1696,n1695);
and gate_1196(n1697,n1691,n1696);
not gate_1197(n1698,n1697);
and gate_1198(n1699,n1531,n1698);
not gate_1199(n1700,n1699);
and gate_1200(n1701,n1677,n1700);
not gate_1201(n1702,n1701);
and gate_1202(n1703,n566,n1702);
not gate_1203(n1704,n1703);
and gate_1204(n1705,pi194,n1701);
not gate_1205(n1706,n1705);
and gate_1206(n1707,n1704,n1706);
not gate_1207(n1708,n1707);
and gate_1208(n1709,n629,n1708);
not gate_1209(n1710,n1709);
and gate_1210(n1711,pi073,n570);
not gate_1211(n1712,n1711);
and gate_1212(n1713,n1710,n1712);
not gate_1213(po062,n1713);
and gate_1214(n1715,pi162,n629);
not gate_1215(n1716,n1715);
and gate_1216(n1717,pi074,n570);
not gate_1217(n1718,n1717);
and gate_1218(n1719,n1716,n1718);
not gate_1219(po063,n1719);
and gate_1220(n1721,n1549,n1602);
not gate_1221(n1722,n1721);
and gate_1222(n1723,n1550,n1574);
not gate_1223(n1724,n1723);
and gate_1224(n1725,n1722,n1724);
not gate_1225(n1726,n1725);
and gate_1226(n1727,n1538,n1544);
not gate_1227(n1728,n1727);
and gate_1228(n1729,n1726,n1727);
not gate_1229(n1730,n1729);
and gate_1230(n1731,n1567,n1574);
not gate_1231(n1732,n1731);
and gate_1232(n1733,n1730,n1732);
not gate_1233(n1734,n1733);
and gate_1234(n1735,n1532,n1734);
not gate_1235(n1736,n1735);
and gate_1236(n1737,n1519,n1607);
not gate_1237(n1738,n1737);
and gate_1238(n1739,n1585,n1738);
and gate_1239(n1740,n1561,n1578);
not gate_1240(n1741,n1740);
and gate_1241(n1742,n1739,n1741);
and gate_1242(n1743,n1519,n1591);
not gate_1243(n1744,n1743);
and gate_1244(n1745,n1563,n1744);
and gate_1245(n1746,n1576,n1745);
and gate_1246(n1747,n1742,n1746);
and gate_1247(n1748,n1593,n1601);
and gate_1248(n1749,n1590,n1748);
and gate_1249(n1750,n1520,n1569);
not gate_1250(n1751,n1750);
and gate_1251(n1752,n1520,n1525);
and gate_1252(n1753,n1579,n1752);
not gate_1253(n1754,n1753);
and gate_1254(n1755,n1751,n1754);
and gate_1255(n1756,n1526,n1583);
and gate_1256(n1757,n1520,n1756);
not gate_1257(n1758,n1757);
and gate_1258(n1759,n1611,n1758);
and gate_1259(n1760,n1755,n1759);
and gate_1260(n1761,n1749,n1760);
and gate_1261(n1762,n1747,n1761);
and gate_1262(n1763,n1519,n1653);
not gate_1263(n1764,n1763);
and gate_1264(n1765,n1525,n1622);
and gate_1265(n1766,n1519,n1765);
not gate_1266(n1767,n1766);
and gate_1267(n1768,n1629,n1767);
and gate_1268(n1769,n1764,n1768);
and gate_1269(n1770,n1519,n1668);
not gate_1270(n1771,n1770);
and gate_1271(n1772,n1624,n1771);
and gate_1272(n1773,n1639,n1772);
and gate_1273(n1774,n1769,n1773);
and gate_1274(n1775,n1520,n1646);
not gate_1275(n1776,n1775);
and gate_1276(n1777,n1670,n1776);
and gate_1277(n1778,n1552,n1603);
not gate_1278(n1779,n1778);
and gate_1279(n1780,n1532,n1644);
and gate_1280(n1781,n1602,n1780);
not gate_1281(n1782,n1781);
and gate_1282(n1783,n1779,n1782);
and gate_1283(n1784,n1777,n1783);
and gate_1284(n1785,n1520,n1765);
not gate_1285(n1786,n1785);
and gate_1286(n1787,n1664,n1786);
and gate_1287(n1788,n1661,n1787);
and gate_1288(n1789,n1784,n1788);
and gate_1289(n1790,n1774,n1789);
and gate_1290(n1791,n1762,n1790);
and gate_1291(n1792,n1736,n1791);
not gate_1292(n1793,n1792);
and gate_1293(n1794,n541,n1793);
not gate_1294(n1795,n1794);
and gate_1295(n1796,pi169,n1792);
not gate_1296(n1797,n1796);
and gate_1297(n1798,n1795,n1797);
not gate_1298(n1799,n1798);
and gate_1299(n1800,n629,n1799);
not gate_1300(n1801,n1800);
and gate_1301(n1802,pi075,n570);
not gate_1302(n1803,n1802);
and gate_1303(n1804,pi067,pi198);
not gate_1304(n1805,n1804);
and gate_1305(n1806,n1803,n1805);
not gate_1306(n1807,n1806);
and gate_1307(n1808,n630,n1807);
not gate_1308(n1809,n1808);
and gate_1309(n1810,n1801,n1809);
not gate_1310(po064,n1810);
and gate_1311(n1812,pi137,n629);
not gate_1312(n1813,n1812);
and gate_1313(n1814,pi076,n570);
not gate_1314(n1815,n1814);
and gate_1315(n1816,pi068,pi198);
not gate_1316(n1817,n1816);
and gate_1317(n1818,n1815,n1817);
not gate_1318(n1819,n1818);
and gate_1319(n1820,n630,n1819);
not gate_1320(n1821,n1820);
and gate_1321(n1822,n1813,n1821);
not gate_1322(po065,n1822);
and gate_1323(n1824,pi157,n581);
not gate_1324(n1825,n1824);
and gate_1325(n1826,n529,pi212);
not gate_1326(n1827,n1826);
and gate_1327(n1828,n1825,n1827);
not gate_1328(n1829,n1828);
and gate_1329(n1830,pi155,n576);
not gate_1330(n1831,n1830);
and gate_1331(n1832,n527,pi206);
not gate_1332(n1833,n1832);
and gate_1333(n1834,n1831,n1833);
not gate_1334(n1835,n1834);
and gate_1335(n1836,pi158,n571);
not gate_1336(n1837,n1836);
and gate_1337(n1838,n530,pi199);
not gate_1338(n1839,n1838);
and gate_1339(n1840,n1837,n1839);
not gate_1340(n1841,n1840);
and gate_1341(n1842,pi159,n592);
not gate_1342(n1843,n1842);
and gate_1343(n1844,n531,pi224);
not gate_1344(n1845,n1844);
and gate_1345(n1846,n1843,n1845);
not gate_1346(n1847,n1846);
and gate_1347(n1848,pi156,n589);
not gate_1348(n1849,n1848);
and gate_1349(n1850,n528,pi221);
not gate_1350(n1851,n1850);
and gate_1351(n1852,n1849,n1851);
not gate_1352(n1853,n1852);
and gate_1353(n1854,n1847,n1853);
not gate_1354(n1855,n1854);
and gate_1355(n1856,n1846,n1852);
not gate_1356(n1857,n1856);
and gate_1357(n1858,n1855,n1857);
not gate_1358(n1859,n1858);
and gate_1359(n1860,n1840,n1859);
and gate_1360(n1861,pi154,n586);
not gate_1361(n1862,n1861);
and gate_1362(n1863,n526,pi217);
not gate_1363(n1864,n1863);
and gate_1364(n1865,n1862,n1864);
not gate_1365(n1866,n1865);
and gate_1366(n1867,n1847,n1865);
not gate_1367(n1868,n1867);
and gate_1368(n1869,n1846,n1866);
not gate_1369(n1870,n1869);
and gate_1370(n1871,n1868,n1870);
and gate_1371(n1872,n1860,n1871);
and gate_1372(n1873,n1835,n1872);
not gate_1373(n1874,n1873);
and gate_1374(n1875,n1841,n1853);
and gate_1375(n1876,n1834,n1869);
and gate_1376(n1877,n1875,n1876);
not gate_1377(n1878,n1877);
and gate_1378(n1879,n1874,n1878);
not gate_1379(n1880,n1879);
and gate_1380(n1881,n1828,n1880);
not gate_1381(n1882,n1881);
and gate_1382(n1883,n1835,n1867);
and gate_1383(n1884,n1840,n1883);
and gate_1384(n1885,n1828,n1884);
and gate_1385(n1886,n1853,n1885);
not gate_1386(n1887,n1886);
and gate_1387(n1888,n1834,n1865);
and gate_1388(n1889,n1847,n1888);
and gate_1389(n1890,n1840,n1889);
and gate_1390(n1891,n1829,n1890);
not gate_1391(n1892,n1891);
and gate_1392(n1893,n1853,n1891);
not gate_1393(n1894,n1893);
and gate_1394(n1895,n1841,n1889);
and gate_1395(n1896,n1828,n1895);
not gate_1396(n1897,n1896);
and gate_1397(n1898,n1852,n1896);
not gate_1398(n1899,n1898);
and gate_1399(n1900,n1894,n1899);
and gate_1400(n1901,n1887,n1900);
and gate_1401(n1902,n1829,n1895);
and gate_1402(n1903,n1852,n1902);
not gate_1403(n1904,n1903);
and gate_1404(n1905,n1841,n1883);
and gate_1405(n1906,n1829,n1905);
not gate_1406(n1907,n1906);
and gate_1407(n1908,n1852,n1906);
not gate_1408(n1909,n1908);
and gate_1409(n1910,n1904,n1909);
and gate_1410(n1911,n1853,n1906);
not gate_1411(n1912,n1911);
and gate_1412(n1913,n1834,n1866);
and gate_1413(n1914,n1847,n1913);
and gate_1414(n1915,n1840,n1914);
and gate_1415(n1916,n1828,n1915);
and gate_1416(n1917,n1852,n1916);
not gate_1417(n1918,n1917);
and gate_1418(n1919,n1912,n1918);
and gate_1419(n1920,n1910,n1919);
and gate_1420(n1921,n1901,n1920);
and gate_1421(n1922,n1829,n1915);
and gate_1422(n1923,n1852,n1922);
not gate_1423(n1924,n1923);
and gate_1424(n1925,n1835,n1866);
and gate_1425(n1926,n1847,n1925);
and gate_1426(n1927,n1840,n1926);
and gate_1427(n1928,n1829,n1927);
and gate_1428(n1929,n1852,n1928);
not gate_1429(n1930,n1929);
and gate_1430(n1931,n1841,n1914);
and gate_1431(n1932,n1828,n1931);
and gate_1432(n1933,n1852,n1932);
not gate_1433(n1934,n1933);
and gate_1434(n1935,n1930,n1934);
and gate_1435(n1936,n1924,n1935);
and gate_1436(n1937,n1853,n1932);
not gate_1437(n1938,n1937);
and gate_1438(n1939,n1841,n1926);
and gate_1439(n1940,n1829,n1939);
and gate_1440(n1941,n1852,n1940);
not gate_1441(n1942,n1941);
and gate_1442(n1943,n1938,n1942);
and gate_1443(n1944,n1853,n1940);
not gate_1444(n1945,n1944);
and gate_1445(n1946,n1846,n1865);
and gate_1446(n1947,n1834,n1946);
and gate_1447(n1948,n1840,n1947);
and gate_1448(n1949,n1828,n1948);
and gate_1449(n1950,n1852,n1949);
not gate_1450(n1951,n1950);
and gate_1451(n1952,n1945,n1951);
and gate_1452(n1953,n1943,n1952);
and gate_1453(n1954,n1936,n1953);
and gate_1454(n1955,n1921,n1954);
and gate_1455(n1956,n1835,n1946);
and gate_1456(n1957,n1841,n1956);
and gate_1457(n1958,n1828,n1957);
not gate_1458(n1959,n1958);
and gate_1459(n1960,n1841,n1947);
and gate_1460(n1961,n1829,n1960);
not gate_1461(n1962,n1961);
and gate_1462(n1963,n1853,n1961);
not gate_1463(n1964,n1963);
and gate_1464(n1965,n1840,n1876);
and gate_1465(n1966,n1828,n1965);
and gate_1466(n1967,n1852,n1966);
not gate_1467(n1968,n1967);
and gate_1468(n1969,n1964,n1968);
and gate_1469(n1970,n1959,n1969);
and gate_1470(n1971,n1828,n1960);
and gate_1471(n1972,n1852,n1971);
not gate_1472(n1973,n1972);
and gate_1473(n1974,n1840,n1956);
and gate_1474(n1975,n1829,n1974);
and gate_1475(n1976,n1852,n1975);
not gate_1476(n1977,n1976);
and gate_1477(n1978,n1829,n1948);
and gate_1478(n1979,n1853,n1978);
not gate_1479(n1980,n1979);
and gate_1480(n1981,n1977,n1980);
and gate_1481(n1982,n1973,n1981);
and gate_1482(n1983,n1970,n1982);
and gate_1483(n1984,n1846,n1925);
and gate_1484(n1985,n1840,n1984);
and gate_1485(n1986,n1828,n1985);
not gate_1486(n1987,n1986);
and gate_1487(n1988,n1829,n1965);
and gate_1488(n1989,n1852,n1988);
not gate_1489(n1990,n1989);
and gate_1490(n1991,n1841,n1984);
and gate_1491(n1992,n1829,n1991);
and gate_1492(n1993,n1852,n1992);
not gate_1493(n1994,n1993);
and gate_1494(n1995,n1990,n1994);
and gate_1495(n1996,n1987,n1995);
and gate_1496(n1997,n1841,n1876);
and gate_1497(n1998,n1829,n1997);
and gate_1498(n1999,n1853,n1998);
not gate_1499(n2000,n1999);
and gate_1500(n2001,n1853,n1992);
not gate_1501(n2002,n2001);
and gate_1502(n2003,n2000,n2002);
and gate_1503(n2004,n1840,n1853);
and gate_1504(n2005,n1829,n2004);
and gate_1505(n2006,n1883,n2005);
not gate_1506(n2007,n2006);
and gate_1507(n2008,n1828,n1853);
and gate_1508(n2009,n1890,n2008);
not gate_1509(n2010,n2009);
and gate_1510(n2011,n2007,n2010);
and gate_1511(n2012,n2003,n2011);
and gate_1512(n2013,n1996,n2012);
and gate_1513(n2014,n1983,n2013);
and gate_1514(n2015,n1955,n2014);
and gate_1515(n2016,n1882,n2015);
not gate_1516(n2017,n2016);
and gate_1517(n2018,n549,n2017);
not gate_1518(n2019,n2018);
and gate_1519(n2020,pi177,n2016);
not gate_1520(n2021,n2020);
and gate_1521(n2022,n2019,n2021);
not gate_1522(n2023,n2022);
and gate_1523(n2024,n629,n2023);
not gate_1524(n2025,n2024);
and gate_1525(n2026,pi077,n570);
not gate_1526(n2027,n2026);
and gate_1527(n2028,pi069,pi198);
not gate_1528(n2029,n2028);
and gate_1529(n2030,n2027,n2029);
not gate_1530(n2031,n2030);
and gate_1531(n2032,n630,n2031);
not gate_1532(n2033,n2032);
and gate_1533(n2034,n2025,n2033);
not gate_1534(po066,n2034);
and gate_1535(n2036,pi145,n629);
not gate_1536(n2037,n2036);
and gate_1537(n2038,pi078,n570);
not gate_1538(n2039,n2038);
and gate_1539(n2040,pi070,pi198);
not gate_1540(n2041,n2040);
and gate_1541(n2042,n2039,n2041);
not gate_1542(n2043,n2042);
and gate_1543(n2044,n630,n2043);
not gate_1544(n2045,n2044);
and gate_1545(n2046,n2037,n2045);
not gate_1546(po067,n2046);
and gate_1547(n2048,n1560,n1744);
and gate_1548(n2049,n1556,n2048);
and gate_1549(n2050,n1519,n1599);
not gate_1550(n2051,n2050);
and gate_1551(n2052,n1738,n2051);
and gate_1552(n2053,n1586,n2052);
and gate_1553(n2054,n2049,n2053);
and gate_1554(n2055,n1605,n1609);
and gate_1555(n2056,n1754,n1758);
and gate_1556(n2057,n2055,n2056);
and gate_1557(n2058,n1598,n1752);
not gate_1558(n2059,n2058);
and gate_1559(n2060,n1748,n2059);
and gate_1560(n2061,n2057,n2060);
and gate_1561(n2062,n2054,n2061);
and gate_1562(n2063,n1519,n1656);
not gate_1563(n2064,n2063);
and gate_1564(n2065,n1624,n2064);
and gate_1565(n2066,n1764,n2065);
and gate_1566(n2067,n1621,n1636);
and gate_1567(n2068,n1643,n1771);
and gate_1568(n2069,n2067,n2068);
and gate_1569(n2070,n2066,n2069);
and gate_1570(n2071,n1602,n1627);
not gate_1571(n2072,n2071);
and gate_1572(n2073,n1658,n2072);
and gate_1573(n2074,n1655,n2073);
and gate_1574(n2075,n1670,n1786);
and gate_1575(n2076,n1672,n1782);
and gate_1576(n2077,n2075,n2076);
and gate_1577(n2078,n2074,n2077);
and gate_1578(n2079,n2070,n2078);
and gate_1579(n2080,n2062,n2079);
and gate_1580(n2081,n1531,n1561);
not gate_1581(n2082,n2081);
and gate_1582(n2083,n1532,n1752);
not gate_1583(n2084,n2083);
and gate_1584(n2085,n2082,n2084);
not gate_1585(n2086,n2085);
and gate_1586(n2087,n1537,n1543);
not gate_1587(n2088,n2087);
and gate_1588(n2089,n1728,n2088);
not gate_1589(n2090,n2089);
and gate_1590(n2091,n2086,n2090);
and gate_1591(n2092,n1550,n2091);
not gate_1592(n2093,n2092);
and gate_1593(n2094,n2080,n2093);
not gate_1594(n2095,n2094);
and gate_1595(n2096,n557,n2095);
not gate_1596(n2097,n2096);
and gate_1597(n2098,pi185,n2094);
not gate_1598(n2099,n2098);
and gate_1599(n2100,n2097,n2099);
not gate_1600(n2101,n2100);
and gate_1601(n2102,n629,n2101);
not gate_1602(n2103,n2102);
and gate_1603(n2104,pi079,n570);
not gate_1604(n2105,n2104);
and gate_1605(n2106,pi071,pi198);
not gate_1606(n2107,n2106);
and gate_1607(n2108,n2105,n2107);
not gate_1608(n2109,n2108);
and gate_1609(n2110,n630,n2109);
not gate_1610(n2111,n2110);
and gate_1611(n2112,n2103,n2111);
not gate_1612(po068,n2112);
and gate_1613(n2114,pi153,n629);
not gate_1614(n2115,n2114);
and gate_1615(n2116,pi080,n570);
not gate_1616(n2117,n2116);
and gate_1617(n2118,pi072,pi198);
not gate_1618(n2119,n2118);
and gate_1619(n2120,n2117,n2119);
not gate_1620(n2121,n2120);
and gate_1621(n2122,n630,n2121);
not gate_1622(n2123,n2122);
and gate_1623(n2124,n2115,n2123);
not gate_1624(po069,n2124);
and gate_1625(n2126,n1860,n1925);
not gate_1626(n2127,n2126);
and gate_1627(n2128,n1875,n1889);
not gate_1628(n2129,n2128);
and gate_1629(n2130,n2127,n2129);
not gate_1630(n2131,n2130);
and gate_1631(n2132,n1829,n2131);
not gate_1632(n2133,n2132);
and gate_1633(n2134,n1852,n1891);
not gate_1634(n2135,n2134);
and gate_1635(n2136,n1905,n2008);
not gate_1636(n2137,n2136);
and gate_1637(n2138,n2135,n2137);
and gate_1638(n2139,n1887,n2138);
and gate_1639(n2140,n1853,n1916);
not gate_1640(n2141,n2140);
and gate_1641(n2142,n1924,n2141);
and gate_1642(n2143,n1907,n2142);
and gate_1643(n2144,n2139,n2143);
and gate_1644(n2145,n1829,n1931);
and gate_1645(n2146,n1853,n2145);
not gate_1646(n2147,n2146);
and gate_1647(n2148,n1938,n2147);
and gate_1648(n2149,n1974,n2008);
not gate_1649(n2150,n2149);
and gate_1650(n2151,n1951,n2150);
and gate_1651(n2152,n2148,n2151);
and gate_1652(n2153,n1828,n1939);
not gate_1653(n2154,n2153);
and gate_1654(n2155,n1852,n2153);
not gate_1655(n2156,n2155);
and gate_1656(n2157,n1935,n2156);
and gate_1657(n2158,n2152,n2157);
and gate_1658(n2159,n2144,n2158);
and gate_1659(n2160,n1852,n1978);
not gate_1660(n2161,n2160);
and gate_1661(n2162,n1981,n2161);
and gate_1662(n2163,n1852,n1958);
not gate_1663(n2164,n2163);
and gate_1664(n2165,n1829,n1957);
and gate_1665(n2166,n1853,n2165);
not gate_1666(n2167,n2166);
and gate_1667(n2168,n2164,n2167);
and gate_1668(n2169,n1853,n1986);
not gate_1669(n2170,n2169);
and gate_1670(n2171,n1968,n2170);
and gate_1671(n2172,n2168,n2171);
and gate_1672(n2173,n2162,n2172);
and gate_1673(n2174,n1984,n2005);
not gate_1674(n2175,n2174);
and gate_1675(n2176,n1990,n2175);
and gate_1676(n2177,n1852,n1998);
not gate_1677(n2178,n2177);
and gate_1678(n2179,n1991,n2008);
not gate_1679(n2180,n2179);
and gate_1680(n2181,n2178,n2180);
and gate_1681(n2182,n2176,n2181);
and gate_1682(n2183,n1852,n1885);
not gate_1683(n2184,n2183);
and gate_1684(n2185,n2010,n2184);
and gate_1685(n2186,n1960,n2008);
not gate_1686(n2187,n2186);
and gate_1687(n2188,n2000,n2187);
and gate_1688(n2189,n2185,n2188);
and gate_1689(n2190,n2182,n2189);
and gate_1690(n2191,n2173,n2190);
and gate_1691(n2192,n2159,n2191);
and gate_1692(n2193,n2133,n2192);
not gate_1693(n2194,n2193);
and gate_1694(n2195,n565,n2194);
not gate_1695(n2196,n2195);
and gate_1696(n2197,pi193,n2193);
not gate_1697(n2198,n2197);
and gate_1698(n2199,n2196,n2198);
not gate_1699(n2200,n2199);
and gate_1700(n2201,n629,n2200);
not gate_1701(n2202,n2201);
and gate_1702(n2203,pi081,n570);
not gate_1703(n2204,n2203);
and gate_1704(n2205,pi073,pi198);
not gate_1705(n2206,n2205);
and gate_1706(n2207,n2204,n2206);
not gate_1707(n2208,n2207);
and gate_1708(n2209,n630,n2208);
not gate_1709(n2210,n2209);
and gate_1710(n2211,n2202,n2210);
not gate_1711(po070,n2211);
and gate_1712(n2213,pi161,n629);
not gate_1713(n2214,n2213);
and gate_1714(n2215,pi082,n570);
not gate_1715(n2216,n2215);
and gate_1716(n2217,pi074,pi198);
not gate_1717(n2218,n2217);
and gate_1718(n2219,n2216,n2218);
not gate_1719(n2220,n2219);
and gate_1720(n2221,n630,n2220);
not gate_1721(n2222,n2221);
and gate_1722(n2223,n2214,n2222);
not gate_1723(po071,n2223);
and gate_1724(n2225,pi134,n607);
not gate_1725(n2226,n2225);
and gate_1726(n2227,n506,pi241);
not gate_1727(n2228,n2227);
and gate_1728(n2229,n2226,n2228);
not gate_1729(n2230,n2229);
and gate_1730(n2231,pi135,n604);
not gate_1731(n2232,n2231);
and gate_1732(n2233,n507,pi237);
not gate_1733(n2234,n2233);
and gate_1734(n2235,n2232,n2234);
not gate_1735(n2236,n2235);
and gate_1736(n2237,pi131,n618);
not gate_1737(n2238,n2237);
and gate_1738(n2239,n503,pi254);
not gate_1739(n2240,n2239);
and gate_1740(n2241,n2238,n2240);
not gate_1741(n2242,n2241);
and gate_1742(n2243,pi133,n600);
not gate_1743(n2244,n2243);
and gate_1744(n2245,n505,pi233);
not gate_1745(n2246,n2245);
and gate_1746(n2247,n2244,n2246);
not gate_1747(n2248,n2247);
and gate_1748(n2249,pi162,n615);
not gate_1749(n2250,n2249);
and gate_1750(n2251,n534,pi251);
not gate_1751(n2252,n2251);
and gate_1752(n2253,n2250,n2252);
not gate_1753(n2254,n2253);
and gate_1754(n2255,n2248,n2254);
not gate_1755(n2256,n2255);
and gate_1756(n2257,n2247,n2253);
not gate_1757(n2258,n2257);
and gate_1758(n2259,n2256,n2258);
not gate_1759(n2260,n2259);
and gate_1760(n2261,pi132,n612);
not gate_1761(n2262,n2261);
and gate_1762(n2263,n504,pi247);
not gate_1763(n2264,n2263);
and gate_1764(n2265,n2262,n2264);
not gate_1765(n2266,n2265);
and gate_1766(n2267,n2254,n2265);
not gate_1767(n2268,n2267);
and gate_1768(n2269,n2253,n2266);
not gate_1769(n2270,n2269);
and gate_1770(n2271,n2268,n2270);
not gate_1771(n2272,n2271);
and gate_1772(n2273,n2260,n2272);
and gate_1773(n2274,n2241,n2273);
and gate_1774(n2275,n2236,n2274);
not gate_1775(n2276,n2275);
and gate_1776(n2277,n2242,n2260);
and gate_1777(n2278,n2266,n2277);
and gate_1778(n2279,n2235,n2278);
not gate_1779(n2280,n2279);
and gate_1780(n2281,n2276,n2280);
not gate_1781(n2282,n2281);
and gate_1782(n2283,n2229,n2282);
not gate_1783(n2284,n2283);
and gate_1784(n2285,n2229,n2235);
and gate_1785(n2286,n2248,n2285);
and gate_1786(n2287,n2265,n2286);
and gate_1787(n2288,n2241,n2287);
and gate_1788(n2289,n2253,n2288);
not gate_1789(n2290,n2289);
and gate_1790(n2291,n2242,n2287);
and gate_1791(n2292,n2253,n2291);
not gate_1792(n2293,n2292);
and gate_1793(n2294,n2290,n2293);
and gate_1794(n2295,n2247,n2285);
and gate_1795(n2296,n2265,n2295);
and gate_1796(n2297,n2241,n2253);
not gate_1797(n2298,n2297);
and gate_1798(n2299,n2296,n2297);
not gate_1799(n2300,n2299);
and gate_1800(n2301,n2294,n2300);
and gate_1801(n2302,n2230,n2235);
and gate_1802(n2303,n2248,n2302);
and gate_1803(n2304,n2265,n2303);
and gate_1804(n2305,n2297,n2304);
not gate_1805(n2306,n2305);
and gate_1806(n2307,n2266,n2303);
and gate_1807(n2308,n2242,n2253);
and gate_1808(n2309,n2307,n2308);
not gate_1809(n2310,n2309);
and gate_1810(n2311,n2306,n2310);
and gate_1811(n2312,n2247,n2302);
and gate_1812(n2313,n2266,n2312);
and gate_1813(n2314,n2242,n2313);
and gate_1814(n2315,n2253,n2314);
not gate_1815(n2316,n2315);
and gate_1816(n2317,n2241,n2307);
and gate_1817(n2318,n2253,n2317);
not gate_1818(n2319,n2318);
and gate_1819(n2320,n2316,n2319);
and gate_1820(n2321,n2311,n2320);
and gate_1821(n2322,n2301,n2321);
and gate_1822(n2323,n2266,n2286);
and gate_1823(n2324,n2241,n2323);
and gate_1824(n2325,n2254,n2324);
not gate_1825(n2326,n2325);
and gate_1826(n2327,n2266,n2295);
and gate_1827(n2328,n2241,n2254);
not gate_1828(n2329,n2328);
and gate_1829(n2330,n2327,n2328);
not gate_1830(n2331,n2330);
and gate_1831(n2332,n2326,n2331);
and gate_1832(n2333,n2242,n2254);
not gate_1833(n2334,n2333);
and gate_1834(n2335,n2296,n2333);
not gate_1835(n2336,n2335);
and gate_1836(n2337,n2332,n2336);
and gate_1837(n2338,n2265,n2312);
and gate_1838(n2339,n2241,n2338);
and gate_1839(n2340,n2254,n2339);
not gate_1840(n2341,n2340);
and gate_1841(n2342,n2242,n2338);
and gate_1842(n2343,n2254,n2342);
not gate_1843(n2344,n2343);
and gate_1844(n2345,n2341,n2344);
and gate_1845(n2346,n2241,n2313);
and gate_1846(n2347,n2254,n2346);
not gate_1847(n2348,n2347);
and gate_1848(n2349,n2304,n2333);
not gate_1849(n2350,n2349);
and gate_1850(n2351,n2348,n2350);
and gate_1851(n2352,n2345,n2351);
and gate_1852(n2353,n2337,n2352);
and gate_1853(n2354,n2322,n2353);
and gate_1854(n2355,n2229,n2236);
and gate_1855(n2356,n2248,n2355);
and gate_1856(n2357,n2265,n2356);
and gate_1857(n2358,n2242,n2357);
and gate_1858(n2359,n2253,n2358);
not gate_1859(n2360,n2359);
and gate_1860(n2361,n2266,n2356);
and gate_1861(n2362,n2297,n2361);
not gate_1862(n2363,n2362);
and gate_1863(n2364,n2360,n2363);
and gate_1864(n2365,n2247,n2355);
and gate_1865(n2366,n2265,n2365);
and gate_1866(n2367,n2297,n2366);
not gate_1867(n2368,n2367);
and gate_1868(n2369,n2364,n2368);
and gate_1869(n2370,n2230,n2236);
and gate_1870(n2371,n2248,n2370);
and gate_1871(n2372,n2265,n2371);
and gate_1872(n2373,n2241,n2372);
and gate_1873(n2374,n2253,n2373);
not gate_1874(n2375,n2374);
and gate_1875(n2376,n2247,n2370);
and gate_1876(n2377,n2266,n2376);
and gate_1877(n2378,n2308,n2377);
not gate_1878(n2379,n2378);
and gate_1879(n2380,n2375,n2379);
and gate_1880(n2381,n2265,n2376);
and gate_1881(n2382,n2242,n2381);
and gate_1882(n2383,n2253,n2382);
not gate_1883(n2384,n2383);
and gate_1884(n2385,n2266,n2371);
and gate_1885(n2386,n2241,n2385);
and gate_1886(n2387,n2253,n2386);
not gate_1887(n2388,n2387);
and gate_1888(n2389,n2384,n2388);
and gate_1889(n2390,n2380,n2389);
and gate_1890(n2391,n2369,n2390);
and gate_1891(n2392,n2242,n2372);
and gate_1892(n2393,n2254,n2392);
not gate_1893(n2394,n2393);
and gate_1894(n2395,n2254,n2386);
not gate_1895(n2396,n2395);
and gate_1896(n2397,n2394,n2396);
and gate_1897(n2398,n2254,n2381);
not gate_1898(n2399,n2398);
and gate_1899(n2400,n2397,n2399);
and gate_1900(n2401,n2266,n2365);
and gate_1901(n2402,n2328,n2401);
not gate_1902(n2403,n2402);
and gate_1903(n2404,n2333,n2401);
not gate_1904(n2405,n2404);
and gate_1905(n2406,n2403,n2405);
and gate_1906(n2407,n2333,n2361);
not gate_1907(n2408,n2407);
and gate_1908(n2409,n2406,n2408);
and gate_1909(n2410,n2400,n2409);
and gate_1910(n2411,n2391,n2410);
and gate_1911(n2412,n2354,n2411);
and gate_1912(n2413,n2284,n2412);
not gate_1913(n2414,n2413);
and gate_1914(n2415,n540,n2414);
not gate_1915(n2416,n2415);
and gate_1916(n2417,pi168,n2413);
not gate_1917(n2418,n2417);
and gate_1918(n2419,n2416,n2418);
not gate_1919(n2420,n2419);
and gate_1920(n2421,n629,n2420);
not gate_1921(n2422,n2421);
and gate_1922(n2423,pi083,n570);
not gate_1923(n2424,n2423);
and gate_1924(n2425,pi075,pi198);
not gate_1925(n2426,n2425);
and gate_1926(n2427,n2424,n2426);
not gate_1927(n2428,n2427);
and gate_1928(n2429,n630,n2428);
not gate_1929(n2430,n2429);
and gate_1930(n2431,n2422,n2430);
not gate_1931(po072,n2431);
and gate_1932(n2433,pi136,n629);
not gate_1933(n2434,n2433);
and gate_1934(n2435,pi084,n570);
not gate_1935(n2436,n2435);
and gate_1936(n2437,pi076,pi198);
not gate_1937(n2438,n2437);
and gate_1938(n2439,n2436,n2438);
not gate_1939(n2440,n2439);
and gate_1940(n2441,n630,n2440);
not gate_1941(n2442,n2441);
and gate_1942(n2443,n2434,n2442);
not gate_1943(po073,n2443);
and gate_1944(n2445,pi142,n609);
not gate_1945(n2446,n2445);
and gate_1946(n2447,n514,pi243);
not gate_1947(n2448,n2447);
and gate_1948(n2449,n2446,n2448);
not gate_1949(n2450,n2449);
and gate_1950(n2451,pi143,n617);
not gate_1951(n2452,n2451);
and gate_1952(n2453,n515,pi253);
not gate_1953(n2454,n2453);
and gate_1954(n2455,n2452,n2454);
not gate_1955(n2456,n2455);
and gate_1956(n2457,pi141,n599);
not gate_1957(n2458,n2457);
and gate_1958(n2459,n513,pi232);
not gate_1959(n2460,n2459);
and gate_1960(n2461,n2458,n2460);
not gate_1961(n2462,n2461);
and gate_1962(n2463,n2455,n2461);
and gate_1963(n2464,pi140,n605);
not gate_1964(n2465,n2464);
and gate_1965(n2466,n512,pi238);
not gate_1966(n2467,n2466);
and gate_1967(n2468,n2465,n2467);
not gate_1968(n2469,n2468);
and gate_1969(n2470,pi139,n614);
not gate_1970(n2471,n2470);
and gate_1971(n2472,n511,pi250);
not gate_1972(n2473,n2472);
and gate_1973(n2474,n2471,n2473);
not gate_1974(n2475,n2474);
and gate_1975(n2476,pi138,n602);
not gate_1976(n2477,n2476);
and gate_1977(n2478,n510,pi235);
not gate_1978(n2479,n2478);
and gate_1979(n2480,n2477,n2479);
not gate_1980(n2481,n2480);
and gate_1981(n2482,n2475,n2481);
and gate_1982(n2483,n2468,n2482);
and gate_1983(n2484,n2463,n2483);
not gate_1984(n2485,n2484);
and gate_1985(n2486,n2469,n2481);
and gate_1986(n2487,n2461,n2486);
not gate_1987(n2488,n2487);
and gate_1988(n2489,n2468,n2480);
and gate_1989(n2490,n2462,n2489);
not gate_1990(n2491,n2490);
and gate_1991(n2492,n2488,n2491);
not gate_1992(n2493,n2492);
and gate_1993(n2494,n2456,n2474);
not gate_1994(n2495,n2494);
and gate_1995(n2496,n2493,n2494);
not gate_1996(n2497,n2496);
and gate_1997(n2498,n2485,n2497);
not gate_1998(n2499,n2498);
and gate_1999(n2500,n2450,n2499);
not gate_2000(n2501,n2500);
and gate_2001(n2502,n2449,n2455);
and gate_2002(n2503,n2462,n2502);
and gate_2003(n2504,n2468,n2503);
and gate_2004(n2505,n2474,n2504);
and gate_2005(n2506,n2480,n2505);
not gate_2006(n2507,n2506);
and gate_2007(n2508,n2450,n2455);
not gate_2008(n2509,n2508);
and gate_2009(n2510,n2461,n2508);
and gate_2010(n2511,n2468,n2510);
and gate_2011(n2512,n2475,n2480);
and gate_2012(n2513,n2511,n2512);
not gate_2013(n2514,n2513);
and gate_2014(n2515,n2507,n2514);
and gate_2015(n2516,n2461,n2502);
and gate_2016(n2517,n2469,n2516);
and gate_2017(n2518,n2512,n2517);
not gate_2018(n2519,n2518);
and gate_2019(n2520,n2515,n2519);
and gate_2020(n2521,n2462,n2508);
and gate_2021(n2522,n2468,n2521);
and gate_2022(n2523,n2475,n2522);
and gate_2023(n2524,n2480,n2523);
not gate_2024(n2525,n2524);
and gate_2025(n2526,n2469,n2521);
and gate_2026(n2527,n2474,n2526);
and gate_2027(n2528,n2480,n2527);
not gate_2028(n2529,n2528);
and gate_2029(n2530,n2525,n2529);
and gate_2030(n2531,n2469,n2510);
and gate_2031(n2532,n2474,n2531);
and gate_2032(n2533,n2480,n2532);
not gate_2033(n2534,n2533);
and gate_2034(n2535,n2512,n2526);
not gate_2035(n2536,n2535);
and gate_2036(n2537,n2534,n2536);
and gate_2037(n2538,n2530,n2537);
and gate_2038(n2539,n2520,n2538);
and gate_2039(n2540,n2481,n2532);
not gate_2040(n2541,n2540);
and gate_2041(n2542,n2469,n2503);
and gate_2042(n2543,n2482,n2542);
not gate_2043(n2544,n2543);
and gate_2044(n2545,n2541,n2544);
and gate_2045(n2546,n2481,n2523);
not gate_2046(n2547,n2546);
and gate_2047(n2548,n2481,n2527);
not gate_2048(n2549,n2548);
and gate_2049(n2550,n2547,n2549);
and gate_2050(n2551,n2545,n2550);
and gate_2051(n2552,n2474,n2542);
and gate_2052(n2553,n2481,n2552);
not gate_2053(n2554,n2553);
and gate_2054(n2555,n2481,n2505);
not gate_2055(n2556,n2555);
and gate_2056(n2557,n2468,n2516);
and gate_2057(n2558,n2482,n2557);
not gate_2058(n2559,n2558);
and gate_2059(n2560,n2556,n2559);
and gate_2060(n2561,n2554,n2560);
and gate_2061(n2562,n2551,n2561);
and gate_2062(n2563,n2539,n2562);
and gate_2063(n2564,n2449,n2456);
not gate_2064(n2565,n2564);
and gate_2065(n2566,n2461,n2564);
and gate_2066(n2567,n2468,n2566);
and gate_2067(n2568,n2474,n2567);
and gate_2068(n2569,n2480,n2568);
not gate_2069(n2570,n2569);
and gate_2070(n2571,n2469,n2566);
and gate_2071(n2572,n2480,n2571);
not gate_2072(n2573,n2572);
and gate_2073(n2574,n2570,n2573);
and gate_2074(n2575,n2462,n2564);
and gate_2075(n2576,n2469,n2575);
and gate_2076(n2577,n2475,n2576);
and gate_2077(n2578,n2480,n2577);
not gate_2078(n2579,n2578);
and gate_2079(n2580,n2450,n2456);
and gate_2080(n2581,n2461,n2580);
and gate_2081(n2582,n2468,n2581);
and gate_2082(n2583,n2474,n2582);
and gate_2083(n2584,n2480,n2583);
not gate_2084(n2585,n2584);
and gate_2085(n2586,n2579,n2585);
and gate_2086(n2587,n2462,n2580);
and gate_2087(n2588,n2469,n2587);
and gate_2088(n2589,n2474,n2588);
and gate_2089(n2590,n2480,n2589);
not gate_2090(n2591,n2590);
and gate_2091(n2592,n2468,n2587);
and gate_2092(n2593,n2512,n2592);
not gate_2093(n2594,n2593);
and gate_2094(n2595,n2591,n2594);
and gate_2095(n2596,n2586,n2595);
and gate_2096(n2597,n2574,n2596);
and gate_2097(n2598,n2475,n2567);
and gate_2098(n2599,n2481,n2598);
not gate_2099(n2600,n2599);
and gate_2100(n2601,n2468,n2575);
and gate_2101(n2602,n2474,n2481);
and gate_2102(n2603,n2601,n2602);
not gate_2103(n2604,n2603);
and gate_2104(n2605,n2600,n2604);
and gate_2105(n2606,n2474,n2576);
and gate_2106(n2607,n2481,n2606);
not gate_2107(n2608,n2607);
and gate_2108(n2609,n2482,n2601);
not gate_2109(n2610,n2609);
and gate_2110(n2611,n2608,n2610);
and gate_2111(n2612,n2605,n2611);
and gate_2112(n2613,n2481,n2583);
not gate_2113(n2614,n2613);
and gate_2114(n2615,n2469,n2581);
and gate_2115(n2616,n2475,n2615);
and gate_2116(n2617,n2481,n2616);
not gate_2117(n2618,n2617);
and gate_2118(n2619,n2614,n2618);
and gate_2119(n2620,n2475,n2588);
and gate_2120(n2621,n2481,n2620);
not gate_2121(n2622,n2621);
and gate_2122(n2623,n2512,n2557);
not gate_2123(n2624,n2623);
and gate_2124(n2625,n2622,n2624);
and gate_2125(n2626,n2619,n2625);
and gate_2126(n2627,n2612,n2626);
and gate_2127(n2628,n2597,n2627);
and gate_2128(n2629,n2563,n2628);
and gate_2129(n2630,n2501,n2629);
not gate_2130(n2631,n2630);
and gate_2131(n2632,n548,n2631);
not gate_2132(n2633,n2632);
and gate_2133(n2634,pi176,n2630);
not gate_2134(n2635,n2634);
and gate_2135(n2636,n2633,n2635);
not gate_2136(n2637,n2636);
and gate_2137(n2638,n629,n2637);
not gate_2138(n2639,n2638);
and gate_2139(n2640,pi085,n570);
not gate_2140(n2641,n2640);
and gate_2141(n2642,pi077,pi198);
not gate_2142(n2643,n2642);
and gate_2143(n2644,n2641,n2643);
not gate_2144(n2645,n2644);
and gate_2145(n2646,n630,n2645);
not gate_2146(n2647,n2646);
and gate_2147(n2648,n2639,n2647);
not gate_2148(po074,n2648);
and gate_2149(n2650,pi144,n629);
not gate_2150(n2651,n2650);
and gate_2151(n2652,pi086,n570);
not gate_2152(n2653,n2652);
and gate_2153(n2654,pi078,pi198);
not gate_2154(n2655,n2654);
and gate_2155(n2656,n2653,n2655);
not gate_2156(n2657,n2656);
and gate_2157(n2658,n630,n2657);
not gate_2158(n2659,n2658);
and gate_2159(n2660,n2651,n2659);
not gate_2160(po075,n2660);
and gate_2161(n2662,n2474,n2517);
and gate_2162(n2663,n2480,n2662);
not gate_2163(n2664,n2663);
and gate_2164(n2665,n2480,n2552);
not gate_2165(n2666,n2665);
and gate_2166(n2667,n2519,n2666);
and gate_2167(n2668,n2664,n2667);
and gate_2168(n2669,n2474,n2522);
and gate_2169(n2670,n2480,n2669);
not gate_2170(n2671,n2670);
and gate_2171(n2672,n2525,n2671);
and gate_2172(n2673,n2537,n2672);
and gate_2173(n2674,n2668,n2673);
and gate_2174(n2675,n2474,n2557);
and gate_2175(n2676,n2481,n2675);
not gate_2176(n2677,n2676);
and gate_2177(n2678,n2560,n2677);
and gate_2178(n2679,n2511,n2602);
not gate_2179(n2680,n2679);
and gate_2180(n2681,n2482,n2531);
not gate_2181(n2682,n2681);
and gate_2182(n2683,n2680,n2682);
and gate_2183(n2684,n2550,n2683);
and gate_2184(n2685,n2678,n2684);
and gate_2185(n2686,n2674,n2685);
and gate_2186(n2687,n2480,n2616);
not gate_2187(n2688,n2687);
and gate_2188(n2689,n2585,n2688);
and gate_2189(n2690,n2480,n2620);
not gate_2190(n2691,n2690);
and gate_2191(n2692,n2591,n2691);
and gate_2192(n2693,n2689,n2692);
and gate_2193(n2694,n2480,n2598);
not gate_2194(n2695,n2694);
and gate_2195(n2696,n2474,n2572);
not gate_2196(n2697,n2696);
and gate_2197(n2698,n2695,n2697);
and gate_2198(n2699,n2579,n2698);
and gate_2199(n2700,n2693,n2699);
and gate_2200(n2701,n2481,n2577);
not gate_2201(n2702,n2701);
and gate_2202(n2703,n2608,n2702);
and gate_2203(n2704,n2600,n2703);
and gate_2204(n2705,n2482,n2582);
not gate_2205(n2706,n2705);
and gate_2206(n2707,n2618,n2706);
and gate_2207(n2708,n2592,n2602);
not gate_2208(n2709,n2708);
and gate_2209(n2710,n2614,n2709);
and gate_2210(n2711,n2707,n2710);
and gate_2211(n2712,n2704,n2711);
and gate_2212(n2713,n2700,n2712);
and gate_2213(n2714,n2686,n2713);
and gate_2214(n2715,n2455,n2475);
not gate_2215(n2716,n2715);
and gate_2216(n2717,n2495,n2716);
not gate_2217(n2718,n2717);
and gate_2218(n2719,n2493,n2718);
and gate_2219(n2720,n2449,n2719);
not gate_2220(n2721,n2720);
and gate_2221(n2722,n2714,n2721);
not gate_2222(n2723,n2722);
and gate_2223(n2724,n556,n2723);
not gate_2224(n2725,n2724);
and gate_2225(n2726,pi184,n2722);
not gate_2226(n2727,n2726);
and gate_2227(n2728,n2725,n2727);
not gate_2228(n2729,n2728);
and gate_2229(n2730,n629,n2729);
not gate_2230(n2731,n2730);
and gate_2231(n2732,pi087,n570);
not gate_2232(n2733,n2732);
and gate_2233(n2734,pi079,pi198);
not gate_2234(n2735,n2734);
and gate_2235(n2736,n2733,n2735);
not gate_2236(n2737,n2736);
and gate_2237(n2738,n630,n2737);
not gate_2238(n2739,n2738);
and gate_2239(n2740,n2731,n2739);
not gate_2240(po076,n2740);
and gate_2241(n2742,pi152,n629);
not gate_2242(n2743,n2742);
and gate_2243(n2744,pi088,n570);
not gate_2244(n2745,n2744);
and gate_2245(n2746,pi080,pi198);
not gate_2246(n2747,n2746);
and gate_2247(n2748,n2745,n2747);
not gate_2248(n2749,n2748);
and gate_2249(n2750,n630,n2749);
not gate_2250(n2751,n2750);
and gate_2251(n2752,n2743,n2751);
not gate_2252(po077,n2752);
and gate_2253(n2754,n1022,n1040);
not gate_2254(n2755,n2754);
and gate_2255(n2756,n1021,n1039);
not gate_2256(n2757,n2756);
and gate_2257(n2758,n2755,n2757);
not gate_2258(n2759,n2758);
and gate_2259(n2760,n1186,n2759);
and gate_2260(n2761,n1027,n2760);
and gate_2261(n2762,n1046,n2761);
not gate_2262(n2763,n2762);
and gate_2263(n2764,n1028,n2759);
and gate_2264(n2765,n1034,n2764);
and gate_2265(n2766,n1045,n2765);
not gate_2266(n2767,n2766);
and gate_2267(n2768,n2763,n2767);
not gate_2268(n2769,n2768);
and gate_2269(n2770,n1051,n2769);
not gate_2270(n2771,n2770);
and gate_2271(n2772,n1033,n1077);
and gate_2272(n2773,n1068,n2772);
not gate_2273(n2774,n2773);
and gate_2274(n2775,n1062,n2774);
and gate_2275(n2776,n1066,n2775);
and gate_2276(n2777,n1021,n1107);
not gate_2277(n2778,n2777);
and gate_2278(n2779,n1021,n1099);
not gate_2279(n2780,n2779);
and gate_2280(n2781,n2778,n2780);
and gate_2281(n2782,n1080,n2781);
and gate_2282(n2783,n2776,n2782);
and gate_2283(n2784,n1092,n2772);
not gate_2284(n2785,n2784);
and gate_2285(n2786,n1098,n2785);
and gate_2286(n2787,n1022,n1028);
and gate_2287(n2788,n1106,n2787);
not gate_2288(n2789,n2788);
and gate_2289(n2790,n1109,n2789);
and gate_2290(n2791,n2786,n2790);
and gate_2291(n2792,n1022,n1060);
not gate_2292(n2793,n2792);
and gate_2293(n2794,n1091,n2793);
and gate_2294(n2795,n2791,n2794);
and gate_2295(n2796,n2783,n2795);
and gate_2296(n2797,n1021,n1152);
not gate_2297(n2798,n2797);
and gate_2298(n2799,n1126,n2798);
and gate_2299(n2800,n1119,n2799);
and gate_2300(n2801,n1034,n1140);
and gate_2301(n2802,n1028,n2801);
and gate_2302(n2803,n1021,n2802);
not gate_2303(n2804,n2803);
and gate_2304(n2805,n1146,n2804);
and gate_2305(n2806,n1140,n1175);
not gate_2306(n2807,n2806);
and gate_2307(n2808,n2805,n2807);
and gate_2308(n2809,n2800,n2808);
and gate_2309(n2810,n1124,n2787);
not gate_2310(n2811,n2810);
and gate_2311(n2812,n1151,n2811);
and gate_2312(n2813,n1159,n2812);
and gate_2313(n2814,n1028,n1141);
and gate_2314(n2815,n1022,n2814);
not gate_2315(n2816,n2815);
and gate_2316(n2817,n1022,n2802);
not gate_2317(n2818,n2817);
and gate_2318(n2819,n2816,n2818);
and gate_2319(n2820,n1092,n1135);
not gate_2320(n2821,n2820);
and gate_2321(n2822,n1164,n2821);
and gate_2322(n2823,n2819,n2822);
and gate_2323(n2824,n2813,n2823);
and gate_2324(n2825,n2809,n2824);
and gate_2325(n2826,n2796,n2825);
and gate_2326(n2827,n2771,n2826);
not gate_2327(n2828,n2827);
and gate_2328(n2829,n564,n2828);
not gate_2329(n2830,n2829);
and gate_2330(n2831,pi192,n2827);
not gate_2331(n2832,n2831);
and gate_2332(n2833,n2830,n2832);
not gate_2333(n2834,n2833);
and gate_2334(n2835,n629,n2834);
not gate_2335(n2836,n2835);
and gate_2336(n2837,pi089,n570);
not gate_2337(n2838,n2837);
and gate_2338(n2839,pi081,pi198);
not gate_2339(n2840,n2839);
and gate_2340(n2841,n2838,n2840);
not gate_2341(n2842,n2841);
and gate_2342(n2843,n630,n2842);
not gate_2343(n2844,n2843);
and gate_2344(n2845,n2836,n2844);
not gate_2345(po078,n2845);
and gate_2346(n2847,pi160,n629);
not gate_2347(n2848,n2847);
and gate_2348(n2849,pi090,n570);
not gate_2349(n2850,n2849);
and gate_2350(n2851,pi082,pi198);
not gate_2351(n2852,n2851);
and gate_2352(n2853,n2850,n2852);
not gate_2353(n2854,n2853);
and gate_2354(n2855,n630,n2854);
not gate_2355(n2856,n2855);
and gate_2356(n2857,n2848,n2856);
not gate_2357(po079,n2857);
and gate_2358(n2859,n1894,n1897);
and gate_2359(n2860,n1930,n2137);
and gate_2360(n2861,n1919,n2860);
and gate_2361(n2862,n2859,n2861);
and gate_2362(n2863,n1942,n2147);
and gate_2363(n2864,n2151,n2863);
and gate_2364(n2865,n1938,n2154);
and gate_2365(n2866,n2864,n2865);
and gate_2366(n2867,n2862,n2866);
and gate_2367(n2868,n1959,n2161);
and gate_2368(n2869,n1962,n1987);
and gate_2369(n2870,n2868,n2869);
and gate_2370(n2871,n2002,n2178);
and gate_2371(n2872,n2185,n2871);
and gate_2372(n2873,n1828,n1997);
and gate_2373(n2874,n1852,n2873);
not gate_2374(n2875,n2874);
and gate_2375(n2876,n2176,n2875);
and gate_2376(n2877,n2872,n2876);
and gate_2377(n2878,n2870,n2877);
and gate_2378(n2879,n2867,n2878);
and gate_2379(n2880,n1858,n1865);
and gate_2380(n2881,n1835,n2880);
not gate_2381(n2882,n2881);
and gate_2382(n2883,n1854,n1913);
not gate_2383(n2884,n2883);
and gate_2384(n2885,n2882,n2884);
not gate_2385(n2886,n2885);
and gate_2386(n2887,n1829,n2886);
not gate_2387(n2888,n2887);
and gate_2388(n2889,n1876,n2008);
not gate_2389(n2890,n2889);
and gate_2390(n2891,n2888,n2890);
not gate_2391(n2892,n2891);
and gate_2392(n2893,n1840,n2892);
not gate_2393(n2894,n2893);
and gate_2394(n2895,n2879,n2894);
not gate_2395(n2896,n2895);
and gate_2396(n2897,n539,n2896);
not gate_2397(n2898,n2897);
and gate_2398(n2899,pi167,n2895);
not gate_2399(n2900,n2899);
and gate_2400(n2901,n2898,n2900);
not gate_2401(n2902,n2901);
and gate_2402(n2903,n629,n2902);
not gate_2403(n2904,n2903);
and gate_2404(n2905,pi091,n570);
not gate_2405(n2906,n2905);
and gate_2406(n2907,pi083,pi198);
not gate_2407(n2908,n2907);
and gate_2408(n2909,n2906,n2908);
not gate_2409(n2910,n2909);
and gate_2410(n2911,n630,n2910);
not gate_2411(n2912,n2911);
and gate_2412(n2913,n2904,n2912);
not gate_2413(po080,n2913);
and gate_2414(n2915,pi135,n629);
not gate_2415(n2916,n2915);
and gate_2416(n2917,pi092,n570);
not gate_2417(n2918,n2917);
and gate_2418(n2919,pi084,pi198);
not gate_2419(n2920,n2919);
and gate_2420(n2921,n2918,n2920);
not gate_2421(n2922,n2921);
and gate_2422(n2923,n630,n2922);
not gate_2423(n2924,n2923);
and gate_2424(n2925,n2916,n2924);
not gate_2425(po081,n2925);
and gate_2426(n2927,n1556,n1745);
and gate_2427(n2928,n1571,n2051);
and gate_2428(n2929,n1741,n2928);
and gate_2429(n2930,n2927,n2929);
and gate_2430(n2931,n1595,n2059);
and gate_2431(n2932,n1590,n2931);
and gate_2432(n2933,n1606,n1755);
and gate_2433(n2934,n2932,n2933);
and gate_2434(n2935,n2930,n2934);
and gate_2435(n2936,n1621,n1767);
and gate_2436(n2937,n2064,n2936);
and gate_2437(n2938,n1648,n1771);
and gate_2438(n2939,n1639,n2938);
and gate_2439(n2940,n2937,n2939);
and gate_2440(n2941,n1666,n1776);
and gate_2441(n2942,n2076,n2941);
and gate_2442(n2943,n1661,n2072);
and gate_2443(n2944,n2942,n2943);
and gate_2444(n2945,n2940,n2944);
and gate_2445(n2946,n2935,n2945);
and gate_2446(n2947,n1525,n1543);
not gate_2447(n2948,n2947);
and gate_2448(n2949,n1689,n2948);
not gate_2449(n2950,n2949);
and gate_2450(n2951,n1519,n1531);
not gate_2451(n2952,n2951);
and gate_2452(n2953,n2950,n2952);
and gate_2453(n2954,n1532,n1537);
not gate_2454(n2955,n2954);
and gate_2455(n2956,n1679,n2955);
and gate_2456(n2957,n2953,n2956);
and gate_2457(n2958,n1550,n2957);
not gate_2458(n2959,n2958);
and gate_2459(n2960,n2946,n2959);
not gate_2460(n2961,n2960);
and gate_2461(n2962,n547,n2961);
not gate_2462(n2963,n2962);
and gate_2463(n2964,pi175,n2960);
not gate_2464(n2965,n2964);
and gate_2465(n2966,n2963,n2965);
not gate_2466(n2967,n2966);
and gate_2467(n2968,n629,n2967);
not gate_2468(n2969,n2968);
and gate_2469(n2970,pi093,n570);
not gate_2470(n2971,n2970);
and gate_2471(n2972,pi085,pi198);
not gate_2472(n2973,n2972);
and gate_2473(n2974,n2971,n2973);
not gate_2474(n2975,n2974);
and gate_2475(n2976,n630,n2975);
not gate_2476(n2977,n2976);
and gate_2477(n2978,n2969,n2977);
not gate_2478(po082,n2978);
and gate_2479(n2980,pi143,n629);
not gate_2480(n2981,n2980);
and gate_2481(n2982,pi094,n570);
not gate_2482(n2983,n2982);
and gate_2483(n2984,pi086,pi198);
not gate_2484(n2985,n2984);
and gate_2485(n2986,n2983,n2985);
not gate_2486(n2987,n2986);
and gate_2487(n2988,n630,n2987);
not gate_2488(n2989,n2988);
and gate_2489(n2990,n2981,n2989);
not gate_2490(po083,n2990);
and gate_2491(n2992,pi134,n597);
not gate_2492(n2993,n2992);
and gate_2493(n2994,n506,pi230);
not gate_2494(n2995,n2994);
and gate_2495(n2996,n2993,n2995);
not gate_2496(n2997,n2996);
and gate_2497(n2998,pi135,n613);
not gate_2498(n2999,n2998);
and gate_2499(n3000,n507,pi249);
not gate_2500(n3001,n3000);
and gate_2501(n3002,n2999,n3001);
not gate_2502(n3003,n3002);
and gate_2503(n3004,pi136,n595);
not gate_2504(n3005,n3004);
and gate_2505(n3006,n508,pi227);
not gate_2506(n3007,n3006);
and gate_2507(n3008,n3005,n3007);
not gate_2508(n3009,n3008);
and gate_2509(n3010,pi139,n606);
not gate_2510(n3011,n3010);
and gate_2511(n3012,n511,pi239);
not gate_2512(n3013,n3012);
and gate_2513(n3014,n3011,n3013);
not gate_2514(n3015,n3014);
and gate_2515(n3016,pi138,n601);
not gate_2516(n3017,n3016);
and gate_2517(n3018,n510,pi234);
not gate_2518(n3019,n3018);
and gate_2519(n3020,n3017,n3019);
not gate_2520(n3021,n3020);
and gate_2521(n3022,pi137,n610);
not gate_2522(n3023,n3022);
and gate_2523(n3024,n509,pi244);
not gate_2524(n3025,n3024);
and gate_2525(n3026,n3023,n3025);
not gate_2526(n3027,n3026);
and gate_2527(n3028,n3020,n3026);
and gate_2528(n3029,n3014,n3028);
and gate_2529(n3030,n3009,n3029);
and gate_2530(n3031,n3003,n3030);
and gate_2531(n3032,n2996,n3031);
not gate_2532(n3033,n3032);
and gate_2533(n3034,n3014,n3027);
and gate_2534(n3035,n3020,n3034);
and gate_2535(n3036,n3009,n3035);
and gate_2536(n3037,n3003,n3036);
and gate_2537(n3038,n2996,n3037);
not gate_2538(n3039,n3038);
and gate_2539(n3040,n3008,n3035);
and gate_2540(n3041,n2996,n3002);
and gate_2541(n3042,n3040,n3041);
not gate_2542(n3043,n3042);
and gate_2543(n3044,n3039,n3043);
and gate_2544(n3045,n3033,n3044);
and gate_2545(n3046,n3014,n3021);
and gate_2546(n3047,n3026,n3046);
and gate_2547(n3048,n3009,n3047);
and gate_2548(n3049,n3003,n3048);
and gate_2549(n3050,n2996,n3049);
not gate_2550(n3051,n3050);
and gate_2551(n3052,n3021,n3027);
and gate_2552(n3053,n3014,n3052);
and gate_2553(n3054,n3008,n3053);
and gate_2554(n3055,n3041,n3054);
not gate_2555(n3056,n3055);
and gate_2556(n3057,n3051,n3056);
and gate_2557(n3058,n3008,n3047);
and gate_2558(n3059,n3003,n3058);
and gate_2559(n3060,n2996,n3059);
not gate_2560(n3061,n3060);
and gate_2561(n3062,n3009,n3053);
and gate_2562(n3063,n3041,n3062);
not gate_2563(n3064,n3063);
and gate_2564(n3065,n3061,n3064);
and gate_2565(n3066,n3057,n3065);
and gate_2566(n3067,n3045,n3066);
and gate_2567(n3068,n2997,n3031);
not gate_2568(n3069,n3068);
and gate_2569(n3070,n3002,n3058);
and gate_2570(n3071,n2997,n3070);
not gate_2571(n3072,n3071);
and gate_2572(n3073,n3069,n3072);
and gate_2573(n3074,n3008,n3029);
and gate_2574(n3075,n2997,n3002);
and gate_2575(n3076,n3074,n3075);
not gate_2576(n3077,n3076);
and gate_2577(n3078,n3073,n3077);
and gate_2578(n3079,n3002,n3048);
and gate_2579(n3080,n2997,n3079);
not gate_2580(n3081,n3080);
and gate_2581(n3082,n2997,n3049);
not gate_2582(n3083,n3082);
and gate_2583(n3084,n3081,n3083);
and gate_2584(n3085,n3003,n3053);
and gate_2585(n3086,n2997,n3085);
not gate_2586(n3087,n3086);
and gate_2587(n3088,n3084,n3087);
and gate_2588(n3089,n3078,n3088);
and gate_2589(n3090,n3067,n3089);
and gate_2590(n3091,n3015,n3020);
and gate_2591(n3092,n3027,n3091);
and gate_2592(n3093,n3009,n3092);
not gate_2593(n3094,n3093);
and gate_2594(n3095,n3002,n3093);
and gate_2595(n3096,n2996,n3095);
not gate_2596(n3097,n3096);
and gate_2597(n3098,n3026,n3091);
and gate_2598(n3099,n3009,n3098);
and gate_2599(n3100,n2996,n3003);
and gate_2600(n3101,n3099,n3100);
not gate_2601(n3102,n3101);
and gate_2602(n3103,n3008,n3092);
and gate_2603(n3104,n3041,n3103);
not gate_2604(n3105,n3104);
and gate_2605(n3106,n3102,n3105);
and gate_2606(n3107,n3097,n3106);
and gate_2607(n3108,n3015,n3021);
and gate_2608(n3109,n3026,n3108);
and gate_2609(n3110,n3008,n3109);
and gate_2610(n3111,n3003,n3110);
and gate_2611(n3112,n2996,n3111);
not gate_2612(n3113,n3112);
and gate_2613(n3114,n3009,n3109);
and gate_2614(n3115,n3041,n3114);
not gate_2615(n3116,n3115);
and gate_2616(n3117,n3113,n3116);
and gate_2617(n3118,n3003,n3093);
and gate_2618(n3119,n2996,n3118);
not gate_2619(n3120,n3119);
and gate_2620(n3121,n3027,n3108);
and gate_2621(n3122,n3008,n3121);
and gate_2622(n3123,n3100,n3122);
not gate_2623(n3124,n3123);
and gate_2624(n3125,n3120,n3124);
and gate_2625(n3126,n3117,n3125);
and gate_2626(n3127,n3107,n3126);
and gate_2627(n3128,n3002,n3099);
and gate_2628(n3129,n2997,n3128);
not gate_2629(n3130,n3129);
and gate_2630(n3131,n2997,n3118);
not gate_2631(n3132,n3131);
and gate_2632(n3133,n3130,n3132);
and gate_2633(n3134,n3008,n3098);
not gate_2634(n3135,n3134);
and gate_2635(n3136,n3075,n3134);
not gate_2636(n3137,n3136);
and gate_2637(n3138,n3133,n3137);
and gate_2638(n3139,n2997,n3111);
not gate_2639(n3140,n3139);
and gate_2640(n3141,n3003,n3114);
and gate_2641(n3142,n2997,n3141);
not gate_2642(n3143,n3142);
and gate_2643(n3144,n3140,n3143);
and gate_2644(n3145,n3009,n3121);
and gate_2645(n3146,n3003,n3145);
and gate_2646(n3147,n2997,n3146);
not gate_2647(n3148,n3147);
and gate_2648(n3149,n3075,n3122);
not gate_2649(n3150,n3149);
and gate_2650(n3151,n3148,n3150);
and gate_2651(n3152,n3144,n3151);
and gate_2652(n3153,n3138,n3152);
and gate_2653(n3154,n3127,n3153);
and gate_2654(n3155,n3090,n3154);
and gate_2655(n3156,n3003,n3015);
not gate_2656(n3157,n3156);
and gate_2657(n3158,n3002,n3014);
not gate_2658(n3159,n3158);
and gate_2659(n3160,n3157,n3159);
not gate_2660(n3161,n3160);
and gate_2661(n3162,n2997,n3027);
not gate_2662(n3163,n3162);
and gate_2663(n3164,n2996,n3026);
not gate_2664(n3165,n3164);
and gate_2665(n3166,n3163,n3165);
not gate_2666(n3167,n3166);
and gate_2667(n3168,n3008,n3167);
and gate_2668(n3169,n3161,n3168);
and gate_2669(n3170,n3020,n3169);
not gate_2670(n3171,n3170);
and gate_2671(n3172,n3155,n3171);
not gate_2672(n3173,n3172);
and gate_2673(n3174,n555,n3173);
not gate_2674(n3175,n3174);
and gate_2675(n3176,pi183,n3172);
not gate_2676(n3177,n3176);
and gate_2677(n3178,n3175,n3177);
not gate_2678(n3179,n3178);
and gate_2679(n3180,n629,n3179);
not gate_2680(n3181,n3180);
and gate_2681(n3182,pi095,n570);
not gate_2682(n3183,n3182);
and gate_2683(n3184,pi087,pi198);
not gate_2684(n3185,n3184);
and gate_2685(n3186,n3183,n3185);
not gate_2686(n3187,n3186);
and gate_2687(n3188,n630,n3187);
not gate_2688(n3189,n3188);
and gate_2689(n3190,n3181,n3189);
not gate_2690(po084,n3190);
and gate_2691(n3192,pi151,n629);
not gate_2692(n3193,n3192);
and gate_2693(n3194,pi096,n570);
not gate_2694(n3195,n3194);
and gate_2695(n3196,pi088,pi198);
not gate_2696(n3197,n3196);
and gate_2697(n3198,n3195,n3197);
not gate_2698(n3199,n3198);
and gate_2699(n3200,n630,n3199);
not gate_2700(n3201,n3200);
and gate_2701(n3202,n3193,n3201);
not gate_2702(po085,n3202);
and gate_2703(n3204,n2480,n2675);
not gate_2704(n3205,n3204);
and gate_2705(n3206,n2519,n2664);
and gate_2706(n3207,n3205,n3206);
and gate_2707(n3208,n2536,n2671);
and gate_2708(n3209,n2515,n3208);
and gate_2709(n3210,n3207,n3209);
and gate_2710(n3211,n2482,n2504);
not gate_2711(n3212,n3211);
and gate_2712(n3213,n2559,n3212);
and gate_2713(n3214,n2677,n3213);
and gate_2714(n3215,n2541,n2682);
and gate_2715(n3216,n2547,n2554);
and gate_2716(n3217,n3215,n3216);
and gate_2717(n3218,n3214,n3217);
and gate_2718(n3219,n3210,n3218);
and gate_2719(n3220,n2570,n2698);
and gate_2720(n3221,n2480,n2606);
not gate_2721(n3222,n3221);
and gate_2722(n3223,n2688,n3222);
and gate_2723(n3224,n2595,n3223);
and gate_2724(n3225,n3220,n3224);
and gate_2725(n3226,n2604,n2608);
and gate_2726(n3227,n2482,n2571);
not gate_2727(n3228,n3227);
and gate_2728(n3229,n3226,n3228);
and gate_2729(n3230,n2614,n2702);
and gate_2730(n3231,n2622,n2706);
and gate_2731(n3232,n3230,n3231);
and gate_2732(n3233,n3229,n3232);
and gate_2733(n3234,n3225,n3233);
and gate_2734(n3235,n3219,n3234);
and gate_2735(n3236,n2450,n2469);
and gate_2736(n3237,n2602,n3236);
not gate_2737(n3238,n3237);
and gate_2738(n3239,n2449,n2468);
and gate_2739(n3240,n2512,n3239);
not gate_2740(n3241,n3240);
and gate_2741(n3242,n3238,n3241);
not gate_2742(n3243,n3242);
and gate_2743(n3244,n2456,n3243);
not gate_2744(n3245,n3244);
and gate_2745(n3246,n2450,n2481);
not gate_2746(n3247,n3246);
and gate_2747(n3248,n2449,n2480);
not gate_2748(n3249,n3248);
and gate_2749(n3250,n3247,n3249);
not gate_2750(n3251,n3250);
and gate_2751(n3252,n2469,n3251);
and gate_2752(n3253,n2715,n3252);
not gate_2753(n3254,n3253);
and gate_2754(n3255,n3245,n3254);
not gate_2755(n3256,n3255);
and gate_2756(n3257,n2462,n3256);
not gate_2757(n3258,n3257);
and gate_2758(n3259,n3235,n3258);
not gate_2759(n3260,n3259);
and gate_2760(n3261,n563,n3260);
not gate_2761(n3262,n3261);
and gate_2762(n3263,pi191,n3259);
not gate_2763(n3264,n3263);
and gate_2764(n3265,n3262,n3264);
not gate_2765(n3266,n3265);
and gate_2766(n3267,n629,n3266);
not gate_2767(n3268,n3267);
and gate_2768(n3269,pi097,n570);
not gate_2769(n3270,n3269);
and gate_2770(n3271,pi089,pi198);
not gate_2771(n3272,n3271);
and gate_2772(n3273,n3270,n3272);
not gate_2773(n3274,n3273);
and gate_2774(n3275,n630,n3274);
not gate_2775(n3276,n3275);
and gate_2776(n3277,n3268,n3276);
not gate_2777(po086,n3277);
and gate_2778(n3279,pi159,n629);
not gate_2779(n3280,n3279);
and gate_2780(n3281,pi098,n570);
not gate_2781(n3282,n3281);
and gate_2782(n3283,pi090,pi198);
not gate_2783(n3284,n3283);
and gate_2784(n3285,n3282,n3284);
not gate_2785(n3286,n3285);
and gate_2786(n3287,n630,n3286);
not gate_2787(n3288,n3287);
and gate_2788(n3289,n3280,n3288);
not gate_2789(po087,n3289);
and gate_2790(n3291,n2667,n3205);
and gate_2791(n3292,n2514,n2671);
and gate_2792(n3293,n2530,n3292);
and gate_2793(n3294,n3291,n3293);
and gate_2794(n3295,n2560,n3212);
and gate_2795(n3296,n2545,n2683);
and gate_2796(n3297,n3295,n3296);
and gate_2797(n3298,n3294,n3297);
and gate_2798(n3299,n2573,n2695);
and gate_2799(n3300,n2585,n3222);
and gate_2800(n3301,n2594,n2691);
and gate_2801(n3302,n3300,n3301);
and gate_2802(n3303,n3299,n3302);
and gate_2803(n3304,n2611,n3228);
and gate_2804(n3305,n2622,n2709);
and gate_2805(n3306,n2707,n3305);
and gate_2806(n3307,n3304,n3306);
and gate_2807(n3308,n3303,n3307);
and gate_2808(n3309,n3298,n3308);
and gate_2809(n3310,n2468,n2565);
not gate_2810(n3311,n3310);
and gate_2811(n3312,n2469,n2564);
not gate_2812(n3313,n3312);
and gate_2813(n3314,n3311,n3313);
and gate_2814(n3315,n2509,n3250);
and gate_2815(n3316,n3314,n3315);
and gate_2816(n3317,n2474,n3316);
not gate_2817(n3318,n3317);
and gate_2818(n3319,n2469,n2512);
and gate_2819(n3320,n2508,n3319);
not gate_2820(n3321,n3320);
and gate_2821(n3322,n3318,n3321);
not gate_2822(n3323,n3322);
and gate_2823(n3324,n2461,n3323);
not gate_2824(n3325,n3324);
and gate_2825(n3326,n3309,n3325);
not gate_2826(n3327,n3326);
and gate_2827(n3328,n538,n3327);
not gate_2828(n3329,n3328);
and gate_2829(n3330,pi166,n3326);
not gate_2830(n3331,n3330);
and gate_2831(n3332,n3329,n3331);
not gate_2832(n3333,n3332);
and gate_2833(n3334,n629,n3333);
not gate_2834(n3335,n3334);
and gate_2835(n3336,pi099,n570);
not gate_2836(n3337,n3336);
and gate_2837(n3338,pi091,pi198);
not gate_2838(n3339,n3338);
and gate_2839(n3340,n3337,n3339);
not gate_2840(n3341,n3340);
and gate_2841(n3342,n630,n3341);
not gate_2842(n3343,n3342);
and gate_2843(n3344,n3335,n3343);
not gate_2844(po088,n3344);
and gate_2845(n3346,pi134,n629);
not gate_2846(n3347,n3346);
and gate_2847(n3348,pi100,n570);
not gate_2848(n3349,n3348);
and gate_2849(n3350,pi092,pi198);
not gate_2850(n3351,n3350);
and gate_2851(n3352,n3349,n3351);
not gate_2852(n3353,n3352);
and gate_2853(n3354,n630,n3353);
not gate_2854(n3355,n3354);
and gate_2855(n3356,n3347,n3355);
not gate_2856(po089,n3356);
and gate_2857(n3358,n2253,n2324);
not gate_2858(n3359,n3358);
and gate_2859(n3360,n2293,n3359);
and gate_2860(n3361,n2300,n3360);
and gate_2861(n3362,n2253,n2342);
not gate_2862(n3363,n3362);
and gate_2863(n3364,n2253,n2346);
not gate_2864(n3365,n3364);
and gate_2865(n3366,n3363,n3365);
and gate_2866(n3367,n2311,n3366);
and gate_2867(n3368,n3361,n3367);
and gate_2868(n3369,n2254,n2291);
not gate_2869(n3370,n3369);
and gate_2870(n3371,n2331,n3370);
and gate_2871(n3372,n2336,n3371);
and gate_2872(n3373,n2326,n2344);
and gate_2873(n3374,n2254,n2314);
not gate_2874(n3375,n3374);
and gate_2875(n3376,n2254,n2317);
not gate_2876(n3377,n3376);
and gate_2877(n3378,n3375,n3377);
and gate_2878(n3379,n3373,n3378);
and gate_2879(n3380,n3372,n3379);
and gate_2880(n3381,n3368,n3380);
and gate_2881(n3382,n2308,n2366);
not gate_2882(n3383,n3382);
and gate_2883(n3384,n2297,n2357);
not gate_2884(n3385,n3384);
and gate_2885(n3386,n3383,n3385);
and gate_2886(n3387,n2368,n3386);
and gate_2887(n3388,n2253,n2392);
not gate_2888(n3389,n3388);
and gate_2889(n3390,n2388,n3389);
and gate_2890(n3391,n2380,n3390);
and gate_2891(n3392,n3387,n3391);
and gate_2892(n3393,n2328,n2381);
not gate_2893(n3394,n3393);
and gate_2894(n3395,n2408,n3394);
and gate_2895(n3396,n2405,n3395);
and gate_2896(n3397,n2241,n2377);
and gate_2897(n3398,n2254,n3397);
not gate_2898(n3399,n3398);
and gate_2899(n3400,n2333,n2385);
not gate_2900(n3401,n3400);
and gate_2901(n3402,n3399,n3401);
and gate_2902(n3403,n2254,n2373);
not gate_2903(n3404,n3403);
and gate_2904(n3405,n2394,n3404);
and gate_2905(n3406,n3402,n3405);
and gate_2906(n3407,n3396,n3406);
and gate_2907(n3408,n3392,n3407);
and gate_2908(n3409,n3381,n3408);
and gate_2909(n3410,n2235,n2329);
not gate_2910(n3411,n3410);
and gate_2911(n3412,n2236,n2241);
not gate_2912(n3413,n3412);
and gate_2913(n3414,n2272,n3413);
and gate_2914(n3415,n3411,n3414);
and gate_2915(n3416,n2247,n3415);
not gate_2916(n3417,n3416);
and gate_2917(n3418,n2248,n2266);
and gate_2918(n3419,n2308,n3418);
not gate_2919(n3420,n3419);
and gate_2920(n3421,n2235,n3419);
not gate_2921(n3422,n3421);
and gate_2922(n3423,n3417,n3422);
not gate_2923(n3424,n3423);
and gate_2924(n3425,n2229,n3424);
not gate_2925(n3426,n3425);
and gate_2926(n3427,n3409,n3426);
not gate_2927(n3428,n3427);
and gate_2928(n3429,n546,n3428);
not gate_2929(n3430,n3429);
and gate_2930(n3431,pi174,n3427);
not gate_2931(n3432,n3431);
and gate_2932(n3433,n3430,n3432);
not gate_2933(n3434,n3433);
and gate_2934(n3435,n629,n3434);
not gate_2935(n3436,n3435);
and gate_2936(n3437,pi101,n570);
not gate_2937(n3438,n3437);
and gate_2938(n3439,pi093,pi198);
not gate_2939(n3440,n3439);
and gate_2940(n3441,n3438,n3440);
not gate_2941(n3442,n3441);
and gate_2942(n3443,n630,n3442);
not gate_2943(n3444,n3443);
and gate_2944(n3445,n3436,n3444);
not gate_2945(po090,n3445);
and gate_2946(n3447,pi142,n629);
not gate_2947(n3448,n3447);
and gate_2948(n3449,pi102,n570);
not gate_2949(n3450,n3449);
and gate_2950(n3451,pi094,pi198);
not gate_2951(n3452,n3451);
and gate_2952(n3453,n3450,n3452);
not gate_2953(n3454,n3453);
and gate_2954(n3455,n630,n3454);
not gate_2955(n3456,n3455);
and gate_2956(n3457,n3448,n3456);
not gate_2957(po091,n3457);
and gate_2958(n3459,n1841,n1865);
not gate_2959(n3460,n3459);
and gate_2960(n3461,n1840,n1866);
not gate_2961(n3462,n3461);
and gate_2962(n3463,n3460,n3462);
not gate_2963(n3464,n3463);
and gate_2964(n3465,n1852,n3464);
and gate_2965(n3466,n1847,n3465);
and gate_2966(n3467,n1835,n3466);
not gate_2967(n3468,n3467);
and gate_2968(n3469,n1947,n2004);
not gate_2969(n3470,n3469);
and gate_2970(n3471,n3468,n3470);
not gate_2971(n3472,n3471);
and gate_2972(n3473,n1828,n3472);
not gate_2973(n3474,n3473);
and gate_2974(n3475,n1887,n1892);
and gate_2975(n3476,n1853,n1896);
not gate_2976(n3477,n3476);
and gate_2977(n3478,n1904,n3477);
and gate_2978(n3479,n1919,n3478);
and gate_2979(n3480,n3475,n3479);
and gate_2980(n3481,n1935,n2141);
and gate_2981(n3482,n1853,n2153);
not gate_2982(n3483,n3482);
and gate_2983(n3484,n2147,n3483);
and gate_2984(n3485,n1952,n3484);
and gate_2985(n3486,n3481,n3485);
and gate_2986(n3487,n3480,n3486);
and gate_2987(n3488,n1973,n1977);
and gate_2988(n3489,n2150,n3488);
and gate_2989(n3490,n1853,n1958);
not gate_2990(n3491,n3490);
and gate_2991(n3492,n1852,n1961);
not gate_2992(n3493,n3492);
and gate_2993(n3494,n3491,n3493);
and gate_2994(n3495,n1852,n1986);
not gate_2995(n3496,n3495);
and gate_2996(n3497,n2167,n3496);
and gate_2997(n3498,n3494,n3497);
and gate_2998(n3499,n3489,n3498);
and gate_2999(n3500,n1994,n2000);
and gate_3000(n3501,n1876,n2005);
not gate_3001(n3502,n3501);
and gate_3002(n3503,n2184,n3502);
and gate_3003(n3504,n3500,n3503);
and gate_3004(n3505,n2180,n2876);
and gate_3005(n3506,n3504,n3505);
and gate_3006(n3507,n3499,n3506);
and gate_3007(n3508,n3487,n3507);
and gate_3008(n3509,n3474,n3508);
not gate_3009(n3510,n3509);
and gate_3010(n3511,n554,n3510);
not gate_3011(n3512,n3511);
and gate_3012(n3513,pi182,n3509);
not gate_3013(n3514,n3513);
and gate_3014(n3515,n3512,n3514);
not gate_3015(n3516,n3515);
and gate_3016(n3517,n629,n3516);
not gate_3017(n3518,n3517);
and gate_3018(n3519,pi103,n570);
not gate_3019(n3520,n3519);
and gate_3020(n3521,pi095,pi198);
not gate_3021(n3522,n3521);
and gate_3022(n3523,n3520,n3522);
not gate_3023(n3524,n3523);
and gate_3024(n3525,n630,n3524);
not gate_3025(n3526,n3525);
and gate_3026(n3527,n3518,n3526);
not gate_3027(po092,n3527);
and gate_3028(n3529,pi150,n629);
not gate_3029(n3530,n3529);
and gate_3030(n3531,pi104,n570);
not gate_3031(n3532,n3531);
and gate_3032(n3533,pi096,pi198);
not gate_3033(n3534,n3533);
and gate_3034(n3535,n3532,n3534);
not gate_3035(n3536,n3535);
and gate_3036(n3537,n630,n3536);
not gate_3037(n3538,n3537);
and gate_3038(n3539,n3530,n3538);
not gate_3039(po093,n3539);
and gate_3040(n3541,n2253,n2339);
not gate_3041(n3542,n3541);
and gate_3042(n3543,n3363,n3542);
and gate_3043(n3544,n2320,n3543);
and gate_3044(n3545,n3361,n3544);
and gate_3045(n3546,n2254,n2288);
not gate_3046(n3547,n3546);
and gate_3047(n3548,n2331,n3547);
and gate_3048(n3549,n2336,n3548);
and gate_3049(n3550,n2341,n2350);
and gate_3050(n3551,n3378,n3550);
and gate_3051(n3552,n3549,n3551);
and gate_3052(n3553,n3545,n3552);
and gate_3053(n3554,n2253,n3397);
not gate_3054(n3555,n3554);
and gate_3055(n3556,n2363,n3555);
and gate_3056(n3557,n2380,n3556);
and gate_3057(n3558,n2360,n3386);
and gate_3058(n3559,n3557,n3558);
and gate_3059(n3560,n2254,n2358);
not gate_3060(n3561,n3560);
and gate_3061(n3562,n2408,n3561);
and gate_3062(n3563,n2403,n3562);
and gate_3063(n3564,n2399,n3402);
and gate_3064(n3565,n3563,n3564);
and gate_3065(n3566,n3559,n3565);
and gate_3066(n3567,n3553,n3566);
and gate_3067(n3568,n2229,n2328);
not gate_3068(n3569,n3568);
and gate_3069(n3570,n2230,n2308);
not gate_3070(n3571,n3570);
and gate_3071(n3572,n3569,n3571);
not gate_3072(n3573,n3572);
and gate_3073(n3574,n2248,n3573);
and gate_3074(n3575,n2236,n3574);
not gate_3075(n3576,n3575);
and gate_3076(n3577,n2298,n2334);
not gate_3077(n3578,n3577);
and gate_3078(n3579,n2295,n3578);
not gate_3079(n3580,n3579);
and gate_3080(n3581,n3576,n3580);
not gate_3081(n3582,n3581);
and gate_3082(n3583,n2266,n3582);
not gate_3083(n3584,n3583);
and gate_3084(n3585,n3567,n3584);
not gate_3085(n3586,n3585);
and gate_3086(n3587,n562,n3586);
not gate_3087(n3588,n3587);
and gate_3088(n3589,pi190,n3585);
not gate_3089(n3590,n3589);
and gate_3090(n3591,n3588,n3590);
not gate_3091(n3592,n3591);
and gate_3092(n3593,n629,n3592);
not gate_3093(n3594,n3593);
and gate_3094(n3595,pi105,n570);
not gate_3095(n3596,n3595);
and gate_3096(n3597,pi097,pi198);
not gate_3097(n3598,n3597);
and gate_3098(n3599,n3596,n3598);
not gate_3099(n3600,n3599);
and gate_3100(n3601,n630,n3600);
not gate_3101(n3602,n3601);
and gate_3102(n3603,n3594,n3602);
not gate_3103(po094,n3603);
and gate_3104(n3605,pi158,n629);
not gate_3105(n3606,n3605);
and gate_3106(n3607,pi106,n570);
not gate_3107(n3608,n3607);
and gate_3108(n3609,pi098,pi198);
not gate_3109(n3610,n3609);
and gate_3110(n3611,n3608,n3610);
not gate_3111(n3612,n3611);
and gate_3112(n3613,n630,n3612);
not gate_3113(n3614,n3613);
and gate_3114(n3615,n3606,n3614);
not gate_3115(po095,n3615);
and gate_3116(n3617,pi150,n587);
not gate_3117(n3618,n3617);
and gate_3118(n3619,n522,pi219);
not gate_3119(n3620,n3619);
and gate_3120(n3621,n3618,n3620);
not gate_3121(n3622,n3621);
and gate_3122(n3623,pi151,n573);
not gate_3123(n3624,n3623);
and gate_3124(n3625,n523,pi201);
not gate_3125(n3626,n3625);
and gate_3126(n3627,n3624,n3626);
not gate_3127(n3628,n3627);
and gate_3128(n3629,pi152,n591);
not gate_3129(n3630,n3629);
and gate_3130(n3631,n524,pi223);
not gate_3131(n3632,n3631);
and gate_3132(n3633,n3630,n3632);
not gate_3133(n3634,n3633);
and gate_3134(n3635,pi153,n584);
not gate_3135(n3636,n3635);
and gate_3136(n3637,n525,pi215);
not gate_3137(n3638,n3637);
and gate_3138(n3639,n3636,n3638);
not gate_3139(n3640,n3639);
and gate_3140(n3641,pi155,n575);
not gate_3141(n3642,n3641);
and gate_3142(n3643,n527,pi204);
not gate_3143(n3644,n3643);
and gate_3144(n3645,n3642,n3644);
not gate_3145(n3646,n3645);
and gate_3146(n3647,pi154,n578);
not gate_3147(n3648,n3647);
and gate_3148(n3649,n526,pi208);
not gate_3149(n3650,n3649);
and gate_3150(n3651,n3648,n3650);
not gate_3151(n3652,n3651);
and gate_3152(n3653,n3645,n3651);
and gate_3153(n3654,n3639,n3653);
and gate_3154(n3655,n3633,n3654);
and gate_3155(n3656,n3627,n3655);
and gate_3156(n3657,n3621,n3656);
not gate_3157(n3658,n3657);
and gate_3158(n3659,n3634,n3654);
and gate_3159(n3660,n3628,n3659);
and gate_3160(n3661,n3621,n3660);
not gate_3161(n3662,n3661);
and gate_3162(n3663,n3640,n3653);
and gate_3163(n3664,n3633,n3663);
and gate_3164(n3665,n3627,n3664);
and gate_3165(n3666,n3621,n3665);
not gate_3166(n3667,n3666);
and gate_3167(n3668,n3662,n3667);
and gate_3168(n3669,n3658,n3668);
and gate_3169(n3670,n3634,n3663);
and gate_3170(n3671,n3627,n3670);
and gate_3171(n3672,n3621,n3671);
not gate_3172(n3673,n3672);
and gate_3173(n3674,n3621,n3628);
and gate_3174(n3675,n3664,n3674);
not gate_3175(n3676,n3675);
and gate_3176(n3677,n3673,n3676);
and gate_3177(n3678,n3645,n3652);
and gate_3178(n3679,n3639,n3678);
and gate_3179(n3680,n3634,n3679);
and gate_3180(n3681,n3628,n3680);
and gate_3181(n3682,n3621,n3681);
not gate_3182(n3683,n3682);
and gate_3183(n3684,n3640,n3678);
and gate_3184(n3685,n3633,n3684);
and gate_3185(n3686,n3627,n3685);
and gate_3186(n3687,n3621,n3686);
not gate_3187(n3688,n3687);
and gate_3188(n3689,n3683,n3688);
and gate_3189(n3690,n3677,n3689);
and gate_3190(n3691,n3669,n3690);
and gate_3191(n3692,n3628,n3670);
and gate_3192(n3693,n3622,n3692);
not gate_3193(n3694,n3693);
and gate_3194(n3695,n3622,n3681);
not gate_3195(n3696,n3695);
and gate_3196(n3697,n3694,n3696);
and gate_3197(n3698,n3622,n3628);
not gate_3198(n3699,n3698);
and gate_3199(n3700,n3685,n3698);
not gate_3200(n3701,n3700);
and gate_3201(n3702,n3634,n3684);
and gate_3202(n3703,n3622,n3627);
and gate_3203(n3704,n3702,n3703);
not gate_3204(n3705,n3704);
and gate_3205(n3706,n3701,n3705);
and gate_3206(n3707,n3697,n3706);
and gate_3207(n3708,n3622,n3665);
not gate_3208(n3709,n3708);
and gate_3209(n3710,n3622,n3671);
not gate_3210(n3711,n3710);
and gate_3211(n3712,n3655,n3698);
not gate_3212(n3713,n3712);
and gate_3213(n3714,n3711,n3713);
and gate_3214(n3715,n3709,n3714);
and gate_3215(n3716,n3707,n3715);
and gate_3216(n3717,n3691,n3716);
and gate_3217(n3718,n3646,n3652);
and gate_3218(n3719,n3640,n3718);
and gate_3219(n3720,n3633,n3719);
and gate_3220(n3721,n3628,n3720);
and gate_3221(n3722,n3621,n3721);
not gate_3222(n3723,n3722);
and gate_3223(n3724,n3639,n3718);
and gate_3224(n3725,n3633,n3724);
and gate_3225(n3726,n3621,n3627);
not gate_3226(n3727,n3726);
and gate_3227(n3728,n3725,n3726);
not gate_3228(n3729,n3728);
and gate_3229(n3730,n3723,n3729);
and gate_3230(n3731,n3634,n3719);
and gate_3231(n3732,n3628,n3731);
and gate_3232(n3733,n3621,n3732);
not gate_3233(n3734,n3733);
and gate_3234(n3735,n3726,n3731);
not gate_3235(n3736,n3735);
and gate_3236(n3737,n3734,n3736);
and gate_3237(n3738,n3730,n3737);
and gate_3238(n3739,n3646,n3651);
and gate_3239(n3740,n3639,n3739);
and gate_3240(n3741,n3633,n3740);
and gate_3241(n3742,n3628,n3741);
and gate_3242(n3743,n3621,n3742);
not gate_3243(n3744,n3743);
and gate_3244(n3745,n3640,n3739);
and gate_3245(n3746,n3633,n3745);
and gate_3246(n3747,n3628,n3746);
and gate_3247(n3748,n3621,n3747);
not gate_3248(n3749,n3748);
and gate_3249(n3750,n3744,n3749);
and gate_3250(n3751,n3634,n3745);
and gate_3251(n3752,n3726,n3751);
not gate_3252(n3753,n3752);
and gate_3253(n3754,n3750,n3753);
and gate_3254(n3755,n3738,n3754);
and gate_3255(n3756,n3622,n3742);
not gate_3256(n3757,n3756);
and gate_3257(n3758,n3703,n3746);
not gate_3258(n3759,n3758);
and gate_3259(n3760,n3698,n3751);
not gate_3260(n3761,n3760);
and gate_3261(n3762,n3759,n3761);
and gate_3262(n3763,n3757,n3762);
and gate_3263(n3764,n3698,n3725);
not gate_3264(n3765,n3764);
and gate_3265(n3766,n3634,n3724);
and gate_3266(n3767,n3703,n3766);
not gate_3267(n3768,n3767);
and gate_3268(n3769,n3765,n3768);
and gate_3269(n3770,n3628,n3766);
and gate_3270(n3771,n3622,n3770);
not gate_3271(n3772,n3771);
and gate_3272(n3773,n3627,n3720);
and gate_3273(n3774,n3622,n3773);
not gate_3274(n3775,n3774);
and gate_3275(n3776,n3772,n3775);
and gate_3276(n3777,n3769,n3776);
and gate_3277(n3778,n3763,n3777);
and gate_3278(n3779,n3755,n3778);
and gate_3279(n3780,n3717,n3779);
and gate_3280(n3781,n3639,n3645);
not gate_3281(n3782,n3781);
and gate_3282(n3783,n3621,n3782);
not gate_3283(n3784,n3783);
and gate_3284(n3785,n3640,n3646);
not gate_3285(n3786,n3785);
and gate_3286(n3787,n3784,n3785);
not gate_3287(n3788,n3787);
and gate_3288(n3789,n3783,n3786);
not gate_3289(n3790,n3789);
and gate_3290(n3791,n3788,n3790);
not gate_3291(n3792,n3791);
and gate_3292(n3793,n3634,n3792);
not gate_3293(n3794,n3793);
and gate_3294(n3795,n3622,n3633);
not gate_3295(n3796,n3795);
and gate_3296(n3797,n3781,n3795);
not gate_3297(n3798,n3797);
and gate_3298(n3799,n3794,n3798);
not gate_3299(n3800,n3799);
and gate_3300(n3801,n3627,n3800);
and gate_3301(n3802,n3652,n3801);
not gate_3302(n3803,n3802);
and gate_3303(n3804,n3780,n3803);
not gate_3304(n3805,n3804);
and gate_3305(n3806,n537,n3805);
not gate_3306(n3807,n3806);
and gate_3307(n3808,pi165,n3804);
not gate_3308(n3809,n3808);
and gate_3309(n3810,n3807,n3809);
not gate_3310(n3811,n3810);
and gate_3311(n3812,n629,n3811);
not gate_3312(n3813,n3812);
and gate_3313(n3814,pi107,n570);
not gate_3314(n3815,n3814);
and gate_3315(n3816,pi099,pi198);
not gate_3316(n3817,n3816);
and gate_3317(n3818,n3815,n3817);
not gate_3318(n3819,n3818);
and gate_3319(n3820,n630,n3819);
not gate_3320(n3821,n3820);
and gate_3321(n3822,n3813,n3821);
not gate_3322(po096,n3822);
and gate_3323(n3824,pi133,n629);
not gate_3324(n3825,n3824);
and gate_3325(n3826,pi108,n570);
not gate_3326(n3827,n3826);
and gate_3327(n3828,pi100,pi198);
not gate_3328(n3829,n3828);
and gate_3329(n3830,n3827,n3829);
not gate_3330(n3831,n3830);
and gate_3331(n3832,n630,n3831);
not gate_3332(n3833,n3832);
and gate_3333(n3834,n3825,n3833);
not gate_3334(po097,n3834);
and gate_3335(n3836,n3033,n3043);
and gate_3336(n3837,n3074,n3100);
not gate_3337(n3838,n3837);
and gate_3338(n3839,n3836,n3838);
and gate_3339(n3840,n2996,n3070);
not gate_3340(n3841,n3840);
and gate_3341(n3842,n3051,n3841);
and gate_3342(n3843,n3003,n3054);
and gate_3343(n3844,n2996,n3843);
not gate_3344(n3845,n3844);
and gate_3345(n3846,n3064,n3845);
and gate_3346(n3847,n3842,n3846);
and gate_3347(n3848,n3839,n3847);
and gate_3348(n3849,n2997,n3059);
not gate_3349(n3850,n3849);
and gate_3350(n3851,n3072,n3850);
and gate_3351(n3852,n3087,n3851);
and gate_3352(n3853,n2997,n3037);
not gate_3353(n3854,n3853);
and gate_3354(n3855,n3030,n3075);
not gate_3355(n3856,n3855);
and gate_3356(n3857,n3069,n3856);
and gate_3357(n3858,n3854,n3857);
and gate_3358(n3859,n3852,n3858);
and gate_3359(n3860,n3848,n3859);
and gate_3360(n3861,n2996,n3128);
not gate_3361(n3862,n3861);
and gate_3362(n3863,n3100,n3103);
not gate_3363(n3864,n3863);
and gate_3364(n3865,n3097,n3864);
and gate_3365(n3866,n3862,n3865);
and gate_3366(n3867,n3002,n3110);
and gate_3367(n3868,n2996,n3867);
not gate_3368(n3869,n3868);
and gate_3369(n3870,n3120,n3869);
and gate_3370(n3871,n3117,n3870);
and gate_3371(n3872,n3866,n3871);
and gate_3372(n3873,n3143,n3150);
and gate_3373(n3874,n3002,n3145);
and gate_3374(n3875,n2997,n3874);
not gate_3375(n3876,n3875);
and gate_3376(n3877,n3030,n3041);
not gate_3377(n3878,n3877);
and gate_3378(n3879,n3876,n3878);
and gate_3379(n3880,n3873,n3879);
and gate_3380(n3881,n3094,n3135);
not gate_3381(n3882,n3881);
and gate_3382(n3883,n2997,n3882);
not gate_3383(n3884,n3883);
and gate_3384(n3885,n3880,n3884);
and gate_3385(n3886,n3872,n3885);
and gate_3386(n3887,n3860,n3886);
and gate_3387(n3888,n3008,n3014);
and gate_3388(n3889,n3075,n3888);
not gate_3389(n3890,n3889);
and gate_3390(n3891,n2997,n3009);
not gate_3391(n3892,n3891);
and gate_3392(n3893,n2996,n3008);
not gate_3393(n3894,n3893);
and gate_3394(n3895,n3892,n3894);
and gate_3395(n3896,n3156,n3895);
not gate_3396(n3897,n3896);
and gate_3397(n3898,n3890,n3897);
not gate_3398(n3899,n3898);
and gate_3399(n3900,n3052,n3899);
not gate_3400(n3901,n3900);
and gate_3401(n3902,n3887,n3901);
not gate_3402(n3903,n3902);
and gate_3403(n3904,n545,n3903);
not gate_3404(n3905,n3904);
and gate_3405(n3906,pi173,n3902);
not gate_3406(n3907,n3906);
and gate_3407(n3908,n3905,n3907);
not gate_3408(n3909,n3908);
and gate_3409(n3910,n629,n3909);
not gate_3410(n3911,n3910);
and gate_3411(n3912,pi109,n570);
not gate_3412(n3913,n3912);
and gate_3413(n3914,pi101,pi198);
not gate_3414(n3915,n3914);
and gate_3415(n3916,n3913,n3915);
not gate_3416(n3917,n3916);
and gate_3417(n3918,n630,n3917);
not gate_3418(n3919,n3918);
and gate_3419(n3920,n3911,n3919);
not gate_3420(po098,n3920);
and gate_3421(n3922,pi141,n629);
not gate_3422(n3923,n3922);
and gate_3423(n3924,pi110,n570);
not gate_3424(n3925,n3924);
and gate_3425(n3926,pi102,pi198);
not gate_3426(n3927,n3926);
and gate_3427(n3928,n3925,n3927);
not gate_3428(n3929,n3928);
and gate_3429(n3930,n630,n3929);
not gate_3430(n3931,n3930);
and gate_3431(n3932,n3923,n3931);
not gate_3432(po099,n3932);
and gate_3433(n3934,n1021,n1086);
not gate_3434(n3935,n3934);
and gate_3435(n3936,n1066,n1070);
and gate_3436(n3937,n3935,n3936);
and gate_3437(n3938,n1021,n1103);
not gate_3438(n3939,n3938);
and gate_3439(n3940,n2778,n3939);
and gate_3440(n3941,n1075,n2774);
and gate_3441(n3942,n3940,n3941);
and gate_3442(n3943,n3937,n3942);
and gate_3443(n3944,n1028,n1084);
and gate_3444(n3945,n1184,n3944);
not gate_3445(n3946,n3945);
and gate_3446(n3947,n1090,n3946);
and gate_3447(n3948,n1094,n3947);
and gate_3448(n3949,n2785,n2793);
and gate_3449(n3950,n1102,n3949);
and gate_3450(n3951,n3948,n3950);
and gate_3451(n3952,n3943,n3951);
and gate_3452(n3953,n1064,n2801);
not gate_3453(n3954,n3953);
and gate_3454(n3955,n2804,n3954);
and gate_3455(n3956,n1139,n3955);
and gate_3456(n3957,n1144,n2799);
and gate_3457(n3958,n3956,n3957);
and gate_3458(n3959,n1034,n1064);
and gate_3459(n3960,n1084,n3959);
not gate_3460(n3961,n3960);
and gate_3461(n3962,n2821,n3961);
and gate_3462(n3963,n1167,n3962);
and gate_3463(n3964,n1092,n1116);
not gate_3464(n3965,n3964);
and gate_3465(n3966,n1154,n3965);
and gate_3466(n3967,n2812,n3966);
and gate_3467(n3968,n3963,n3967);
and gate_3468(n3969,n3958,n3968);
and gate_3469(n3970,n3952,n3969);
and gate_3470(n3971,n1040,n1052);
and gate_3471(n3972,n2787,n3971);
not gate_3472(n3973,n3972);
and gate_3473(n3974,n1064,n1083);
not gate_3474(n3975,n3974);
and gate_3475(n3976,n3973,n3975);
not gate_3476(n3977,n3976);
and gate_3477(n3978,n1046,n3977);
not gate_3478(n3979,n3978);
and gate_3479(n3980,n1053,n1172);
not gate_3480(n3981,n3980);
and gate_3481(n3982,n3979,n3981);
not gate_3482(n3983,n3982);
and gate_3483(n3984,n1033,n3983);
not gate_3484(n3985,n3984);
and gate_3485(n3986,n3970,n3985);
not gate_3486(n3987,n3986);
and gate_3487(n3988,n553,n3987);
not gate_3488(n3989,n3988);
and gate_3489(n3990,pi181,n3986);
not gate_3490(n3991,n3990);
and gate_3491(n3992,n3989,n3991);
not gate_3492(n3993,n3992);
and gate_3493(n3994,n629,n3993);
not gate_3494(n3995,n3994);
and gate_3495(n3996,pi111,n570);
not gate_3496(n3997,n3996);
and gate_3497(n3998,pi103,pi198);
not gate_3498(n3999,n3998);
and gate_3499(n4000,n3997,n3999);
not gate_3500(n4001,n4000);
and gate_3501(n4002,n630,n4001);
not gate_3502(n4003,n4002);
and gate_3503(n4004,n3995,n4003);
not gate_3504(po100,n4004);
and gate_3505(n4006,pi149,n629);
not gate_3506(n4007,n4006);
and gate_3507(n4008,pi112,n570);
not gate_3508(n4009,n4008);
and gate_3509(n4010,pi104,pi198);
not gate_3510(n4011,n4010);
and gate_3511(n4012,n4009,n4011);
not gate_3512(n4013,n4012);
and gate_3513(n4014,n630,n4013);
not gate_3514(n4015,n4014);
and gate_3515(n4016,n4007,n4015);
not gate_3516(po101,n4016);
and gate_3517(n4018,n3622,n3656);
not gate_3518(n4019,n4018);
and gate_3519(n4020,n3622,n3660);
not gate_3520(n4021,n4020);
and gate_3521(n4022,n3713,n4021);
and gate_3522(n4023,n4019,n4022);
and gate_3523(n4024,n3627,n3680);
and gate_3524(n4025,n3622,n4024);
not gate_3525(n4026,n4025);
and gate_3526(n4027,n3709,n4026);
and gate_3527(n4028,n3706,n4027);
and gate_3528(n4029,n4023,n4028);
and gate_3529(n4030,n3621,n3692);
not gate_3530(n4031,n4030);
and gate_3531(n4032,n3621,n3633);
and gate_3532(n4033,n3628,n3679);
and gate_3533(n4034,n4032,n4033);
not gate_3534(n4035,n4034);
and gate_3535(n4036,n4031,n4035);
and gate_3536(n4037,n3659,n3726);
not gate_3537(n4038,n4037);
and gate_3538(n4039,n4036,n4038);
and gate_3539(n4040,n3690,n4039);
and gate_3540(n4041,n4029,n4040);
and gate_3541(n4042,n3634,n3740);
and gate_3542(n4043,n3674,n4042);
not gate_3543(n4044,n4043);
and gate_3544(n4045,n3749,n4044);
and gate_3545(n4046,n3726,n3741);
not gate_3546(n4047,n4046);
and gate_3547(n4048,n4045,n4047);
and gate_3548(n4049,n3729,n3753);
and gate_3549(n4050,n3621,n3773);
not gate_3550(n4051,n4050);
and gate_3551(n4052,n3734,n4051);
and gate_3552(n4053,n4049,n4052);
and gate_3553(n4054,n4048,n4053);
and gate_3554(n4055,n3622,n3721);
not gate_3555(n4056,n4055);
and gate_3556(n4057,n3698,n3702);
not gate_3557(n4058,n4057);
and gate_3558(n4059,n4056,n4058);
and gate_3559(n4060,n3776,n4059);
and gate_3560(n4061,n3622,n3747);
not gate_3561(n4062,n4061);
and gate_3562(n4063,n3765,n4062);
and gate_3563(n4064,n3703,n4042);
not gate_3564(n4065,n4064);
and gate_3565(n4066,n3761,n4065);
and gate_3566(n4067,n4063,n4066);
and gate_3567(n4068,n4060,n4067);
and gate_3568(n4069,n4054,n4068);
and gate_3569(n4070,n4041,n4069);
and gate_3570(n4071,n3622,n3651);
not gate_3571(n4072,n4071);
and gate_3572(n4073,n3621,n3652);
not gate_3573(n4074,n4073);
and gate_3574(n4075,n4072,n4074);
not gate_3575(n4076,n4075);
and gate_3576(n4077,n3699,n3727);
and gate_3577(n4078,n4076,n4077);
and gate_3578(n4079,n3646,n4078);
not gate_3579(n4080,n4079);
and gate_3580(n4081,n3678,n3726);
not gate_3581(n4082,n4081);
and gate_3582(n4083,n4080,n4082);
not gate_3583(n4084,n4083);
and gate_3584(n4085,n3633,n4084);
and gate_3585(n4086,n3639,n4085);
not gate_3586(n4087,n4086);
and gate_3587(n4088,n4070,n4087);
not gate_3588(n4089,n4088);
and gate_3589(n4090,n561,n4089);
not gate_3590(n4091,n4090);
and gate_3591(n4092,pi189,n4088);
not gate_3592(n4093,n4092);
and gate_3593(n4094,n4091,n4093);
not gate_3594(n4095,n4094);
and gate_3595(n4096,n629,n4095);
not gate_3596(n4097,n4096);
and gate_3597(n4098,pi113,n570);
not gate_3598(n4099,n4098);
and gate_3599(n4100,pi105,pi198);
not gate_3600(n4101,n4100);
and gate_3601(n4102,n4099,n4101);
not gate_3602(n4103,n4102);
and gate_3603(n4104,n630,n4103);
not gate_3604(n4105,n4104);
and gate_3605(n4106,n4097,n4105);
not gate_3606(po102,n4106);
and gate_3607(n4108,pi157,n629);
not gate_3608(n4109,n4108);
and gate_3609(n4110,pi114,n570);
not gate_3610(n4111,n4110);
and gate_3611(n4112,pi106,pi198);
not gate_3612(n4113,n4112);
and gate_3613(n4114,n4111,n4113);
not gate_3614(n4115,n4114);
and gate_3615(n4116,n630,n4115);
not gate_3616(n4117,n4116);
and gate_3617(n4118,n4109,n4117);
not gate_3618(po103,n4118);
and gate_3619(n4120,n1310,n1313);
and gate_3620(n4121,n1439,n4120);
and gate_3621(n4122,n1275,n1302);
not gate_3622(n4123,n4122);
and gate_3623(n4124,n1336,n4123);
and gate_3624(n4125,n1333,n1443);
and gate_3625(n4126,n4124,n4125);
and gate_3626(n4127,n4121,n4126);
and gate_3627(n4128,n1295,n1437);
and gate_3628(n4129,n1426,n4128);
and gate_3629(n4130,n1289,n4129);
and gate_3630(n4131,n4127,n4130);
and gate_3631(n4132,n1220,n1465);
not gate_3632(n4133,n4132);
and gate_3633(n4134,n1344,n4133);
and gate_3634(n4135,n1450,n4134);
and gate_3635(n4136,n1360,n1458);
and gate_3636(n4137,n1354,n4136);
and gate_3637(n4138,n4135,n4137);
and gate_3638(n4139,n1221,n1448);
not gate_3639(n4140,n4139);
and gate_3640(n4141,n1463,n4140);
and gate_3641(n4142,n1362,n4141);
and gate_3642(n4143,n1370,n1375);
and gate_3643(n4144,n1220,n1429);
not gate_3644(n4145,n4144);
and gate_3645(n4146,n1470,n4145);
and gate_3646(n4147,n4143,n4146);
and gate_3647(n4148,n4142,n4147);
and gate_3648(n4149,n4138,n4148);
and gate_3649(n4150,n4131,n4149);
and gate_3650(n4151,n1227,n1386);
and gate_3651(n4152,n1233,n4151);
and gate_3652(n4153,n1244,n4152);
not gate_3653(n4154,n4153);
and gate_3654(n4155,n1233,n1239);
and gate_3655(n4156,n1302,n4155);
not gate_3656(n4157,n4156);
and gate_3657(n4158,n1232,n1238);
and gate_3658(n4159,n1276,n4158);
not gate_3659(n4160,n4159);
and gate_3660(n4161,n4157,n4160);
not gate_3661(n4162,n4161);
and gate_3662(n4163,n1245,n4162);
not gate_3663(n4164,n4163);
and gate_3664(n4165,n4154,n4164);
not gate_3665(n4166,n4165);
and gate_3666(n4167,n1250,n4166);
not gate_3667(n4168,n4167);
and gate_3668(n4169,n4150,n4168);
not gate_3669(n4170,n4169);
and gate_3670(n4171,n536,n4170);
not gate_3671(n4172,n4171);
and gate_3672(n4173,pi164,n4169);
not gate_3673(n4174,n4173);
and gate_3674(n4175,n4172,n4174);
not gate_3675(n4176,n4175);
and gate_3676(n4177,n629,n4176);
not gate_3677(n4178,n4177);
and gate_3678(n4179,pi115,n570);
not gate_3679(n4180,n4179);
and gate_3680(n4181,pi107,pi198);
not gate_3681(n4182,n4181);
and gate_3682(n4183,n4180,n4182);
not gate_3683(n4184,n4183);
and gate_3684(n4185,n630,n4184);
not gate_3685(n4186,n4185);
and gate_3686(n4187,n4178,n4186);
not gate_3687(po104,n4187);
and gate_3688(n4189,pi132,n629);
not gate_3689(n4190,n4189);
and gate_3690(n4191,pi116,n570);
not gate_3691(n4192,n4191);
and gate_3692(n4193,pi108,pi198);
not gate_3693(n4194,n4193);
and gate_3694(n4195,n4192,n4194);
not gate_3695(n4196,n4195);
and gate_3696(n4197,n630,n4196);
not gate_3697(n4198,n4197);
and gate_3698(n4199,n4190,n4198);
not gate_3699(po105,n4199);
and gate_3700(n4201,n1257,n1278);
and gate_3701(n4202,n1268,n4201);
and gate_3702(n4203,n1288,n1432);
and gate_3703(n4204,n4202,n4203);
and gate_3704(n4205,n1437,n4123);
and gate_3705(n4206,n1299,n4205);
and gate_3706(n4207,n1318,n1327);
and gate_3707(n4208,n4125,n4207);
and gate_3708(n4209,n4206,n4208);
and gate_3709(n4210,n4204,n4209);
and gate_3710(n4211,n1353,n1360);
and gate_3711(n4212,n4141,n4211);
and gate_3712(n4213,n1455,n4134);
and gate_3713(n4214,n4212,n4213);
and gate_3714(n4215,n1371,n1467);
and gate_3715(n4216,n1373,n4145);
and gate_3716(n4217,n1473,n4216);
and gate_3717(n4218,n4215,n4217);
and gate_3718(n4219,n4214,n4218);
and gate_3719(n4220,n4210,n4219);
and gate_3720(n4221,n1385,n1479);
and gate_3721(n4222,n1233,n4221);
and gate_3722(n4223,n1245,n4222);
not gate_3723(n4224,n4223);
and gate_3724(n4225,n1232,n1479);
and gate_3725(n4226,n1239,n4225);
and gate_3726(n4227,n1244,n4226);
not gate_3727(n4228,n4227);
and gate_3728(n4229,n4224,n4228);
not gate_3729(n4230,n4229);
and gate_3730(n4231,n1250,n4230);
not gate_3731(n4232,n4231);
and gate_3732(n4233,n4220,n4232);
not gate_3733(n4234,n4233);
and gate_3734(n4235,n544,n4234);
not gate_3735(n4236,n4235);
and gate_3736(n4237,pi172,n4233);
not gate_3737(n4238,n4237);
and gate_3738(n4239,n4236,n4238);
not gate_3739(n4240,n4239);
and gate_3740(n4241,n629,n4240);
not gate_3741(n4242,n4241);
and gate_3742(n4243,pi117,n570);
not gate_3743(n4244,n4243);
and gate_3744(n4245,pi109,pi198);
not gate_3745(n4246,n4245);
and gate_3746(n4247,n4244,n4246);
not gate_3747(n4248,n4247);
and gate_3748(n4249,n630,n4248);
not gate_3749(n4250,n4249);
and gate_3750(n4251,n4242,n4250);
not gate_3751(po106,n4251);
and gate_3752(n4253,pi140,n629);
not gate_3753(n4254,n4253);
and gate_3754(n4255,pi118,n570);
not gate_3755(n4256,n4255);
and gate_3756(n4257,pi110,pi198);
not gate_3757(n4258,n4257);
and gate_3758(n4259,n4256,n4258);
not gate_3759(n4260,n4259);
and gate_3760(n4261,n630,n4260);
not gate_3761(n4262,n4261);
and gate_3762(n4263,n4254,n4262);
not gate_3763(po107,n4263);
and gate_3764(n4265,n2247,n2265);
and gate_3765(n4266,n2328,n4265);
not gate_3766(n4267,n4266);
and gate_3767(n4268,n3420,n4267);
not gate_3768(n4269,n4268);
and gate_3769(n4270,n2236,n4269);
not gate_3770(n4271,n4270);
and gate_3771(n4272,n2235,n2308);
and gate_3772(n4273,n4265,n4272);
not gate_3773(n4274,n4273);
and gate_3774(n4275,n4271,n4274);
not gate_3775(n4276,n4275);
and gate_3776(n4277,n2229,n4276);
not gate_3777(n4278,n4277);
and gate_3778(n4279,n2290,n3360);
and gate_3779(n4280,n3365,n3542);
and gate_3780(n4281,n2310,n2316);
and gate_3781(n4282,n4280,n4281);
and gate_3782(n4283,n4279,n4282);
and gate_3783(n4284,n3370,n3547);
and gate_3784(n4285,n2336,n4284);
and gate_3785(n4286,n2326,n3375);
and gate_3786(n4287,n2351,n4286);
and gate_3787(n4288,n4285,n4287);
and gate_3788(n4289,n4283,n4288);
and gate_3789(n4290,n2363,n3383);
and gate_3790(n4291,n2368,n4290);
and gate_3791(n4292,n2384,n3555);
and gate_3792(n4293,n2375,n3389);
and gate_3793(n4294,n4292,n4293);
and gate_3794(n4295,n4291,n4294);
and gate_3795(n4296,n3394,n3561);
and gate_3796(n4297,n2406,n4296);
and gate_3797(n4298,n2396,n3404);
and gate_3798(n4299,n2307,n2333);
not gate_3799(n4300,n4299);
and gate_3800(n4301,n3401,n4300);
and gate_3801(n4302,n4298,n4301);
and gate_3802(n4303,n4297,n4302);
and gate_3803(n4304,n4295,n4303);
and gate_3804(n4305,n4289,n4304);
and gate_3805(n4306,n4278,n4305);
not gate_3806(n4307,n4306);
and gate_3807(n4308,n552,n4307);
not gate_3808(n4309,n4308);
and gate_3809(n4310,pi180,n4306);
not gate_3810(n4311,n4310);
and gate_3811(n4312,n4309,n4311);
not gate_3812(n4313,n4312);
and gate_3813(n4314,n629,n4313);
not gate_3814(n4315,n4314);
and gate_3815(n4316,pi119,n570);
not gate_3816(n4317,n4316);
and gate_3817(n4318,pi111,pi198);
not gate_3818(n4319,n4318);
and gate_3819(n4320,n4317,n4319);
not gate_3820(n4321,n4320);
and gate_3821(n4322,n630,n4321);
not gate_3822(n4323,n4322);
and gate_3823(n4324,n4315,n4323);
not gate_3824(po108,n4324);
and gate_3825(n4326,pi148,n629);
not gate_3826(n4327,n4326);
and gate_3827(n4328,pi120,n570);
not gate_3828(n4329,n4328);
and gate_3829(n4330,pi112,pi198);
not gate_3830(n4331,n4330);
and gate_3831(n4332,n4329,n4331);
not gate_3832(n4333,n4332);
and gate_3833(n4334,n630,n4333);
not gate_3834(n4335,n4334);
and gate_3835(n4336,n4327,n4335);
not gate_3836(po109,n4336);
and gate_3837(n4338,n3015,n3168);
not gate_3838(n4339,n4338);
and gate_3839(n4340,n3034,n3891);
not gate_3840(n4341,n4340);
and gate_3841(n4342,n4339,n4341);
not gate_3842(n4343,n4342);
and gate_3843(n4344,n3002,n4343);
and gate_3844(n4345,n3020,n4344);
not gate_3845(n4346,n4345);
and gate_3846(n4347,n3044,n3838);
and gate_3847(n4348,n2996,n3079);
not gate_3848(n4349,n4348);
and gate_3849(n4350,n3841,n4349);
and gate_3850(n4351,n3057,n4350);
and gate_3851(n4352,n4347,n4351);
and gate_3852(n4353,n3077,n3857);
and gate_3853(n4354,n3003,n3040);
and gate_3854(n4355,n2997,n4354);
not gate_3855(n4356,n4355);
and gate_3856(n4357,n3850,n4356);
and gate_3857(n4358,n2997,n3843);
not gate_3858(n4359,n4358);
and gate_3859(n4360,n3081,n4359);
and gate_3860(n4361,n4357,n4360);
and gate_3861(n4362,n4353,n4361);
and gate_3862(n4363,n4352,n4362);
and gate_3863(n4364,n3102,n3864);
and gate_3864(n4365,n3862,n4364);
and gate_3865(n4366,n2996,n3874);
not gate_3866(n4367,n4366);
and gate_3867(n4368,n3113,n4367);
and gate_3868(n4369,n3097,n3124);
and gate_3869(n4370,n4368,n4369);
and gate_3870(n4371,n4365,n4370);
and gate_3871(n4372,n3062,n3100);
not gate_3872(n4373,n4372);
and gate_3873(n4374,n3876,n4373);
and gate_3874(n4375,n3144,n4374);
and gate_3875(n4376,n3003,n3134);
and gate_3876(n4377,n2997,n4376);
not gate_3877(n4378,n4377);
and gate_3878(n4379,n2997,n3867);
not gate_3879(n4380,n4379);
and gate_3880(n4381,n4378,n4380);
and gate_3881(n4382,n3133,n4381);
and gate_3882(n4383,n4375,n4382);
and gate_3883(n4384,n4371,n4383);
and gate_3884(n4385,n4363,n4384);
and gate_3885(n4386,n4346,n4385);
not gate_3886(n4387,n4386);
and gate_3887(n4388,n560,n4387);
not gate_3888(n4389,n4388);
and gate_3889(n4390,pi188,n4386);
not gate_3890(n4391,n4390);
and gate_3891(n4392,n4389,n4391);
not gate_3892(n4393,n4392);
and gate_3893(n4394,n629,n4393);
not gate_3894(n4395,n4394);
and gate_3895(n4396,pi113,pi198);
not gate_3896(n4397,n4396);
and gate_3897(n4398,pi121,n570);
not gate_3898(n4399,n4398);
and gate_3899(n4400,n4397,n4399);
not gate_3900(n4401,n4400);
and gate_3901(n4402,n630,n4401);
not gate_3902(n4403,n4402);
and gate_3903(n4404,n4395,n4403);
not gate_3904(po110,n4404);
and gate_3905(n4406,pi156,n629);
not gate_3906(n4407,n4406);
and gate_3907(n4408,pi114,pi198);
not gate_3908(n4409,n4408);
and gate_3909(n4410,pi122,n570);
not gate_3910(n4411,n4410);
and gate_3911(n4412,n4409,n4411);
not gate_3912(n4413,n4412);
and gate_3913(n4414,n630,n4413);
not gate_3914(n4415,n4414);
and gate_3915(n4416,n4407,n4415);
not gate_3916(po111,n4416);
and gate_3917(n4418,n3039,n3061);
and gate_3918(n4419,n3845,n4349);
and gate_3919(n4420,n4418,n4419);
and gate_3920(n4421,n3839,n4420);
and gate_3921(n4422,n3856,n4356);
and gate_3922(n4423,n3077,n4422);
and gate_3923(n4424,n3072,n3854);
and gate_3924(n4425,n3083,n4359);
and gate_3925(n4426,n4424,n4425);
and gate_3926(n4427,n4423,n4426);
and gate_3927(n4428,n4421,n4427);
and gate_3928(n4429,n3106,n3862);
and gate_3929(n4430,n3870,n4368);
and gate_3930(n4431,n4429,n4430);
and gate_3931(n4432,n2997,n3095);
not gate_3932(n4433,n4432);
and gate_3933(n4434,n3130,n4433);
and gate_3934(n4435,n4378,n4434);
and gate_3935(n4436,n3143,n4380);
and gate_3936(n4437,n3151,n4436);
and gate_3937(n4438,n4435,n4437);
and gate_3938(n4439,n4431,n4438);
and gate_3939(n4440,n4428,n4439);
and gate_3940(n4441,n2997,n3021);
not gate_3941(n4442,n4441);
and gate_3942(n4443,n2996,n3020);
not gate_3943(n4444,n4443);
and gate_3944(n4445,n4442,n4444);
not gate_3945(n4446,n4445);
and gate_3946(n4447,n3026,n4445);
and gate_3947(n4448,n3156,n4447);
not gate_3948(n4449,n4448);
and gate_3949(n4450,n3002,n4446);
and gate_3950(n4451,n3034,n4450);
not gate_3951(n4452,n4451);
and gate_3952(n4453,n4449,n4452);
not gate_3953(n4454,n4453);
and gate_3954(n4455,n3009,n4454);
not gate_3955(n4456,n4455);
and gate_3956(n4457,n4440,n4456);
not gate_3957(n4458,n4457);
and gate_3958(n4459,n535,n4458);
not gate_3959(n4460,n4459);
and gate_3960(n4461,pi163,n4457);
not gate_3961(n4462,n4461);
and gate_3962(n4463,n4460,n4462);
not gate_3963(n4464,n4463);
and gate_3964(n4465,n629,n4464);
not gate_3965(n4466,n4465);
and gate_3966(n4467,pi115,pi198);
not gate_3967(n4468,n4467);
and gate_3968(n4469,pi123,n570);
not gate_3969(n4470,n4469);
and gate_3970(n4471,n4468,n4470);
not gate_3971(n4472,n4471);
and gate_3972(n4473,n630,n4472);
not gate_3973(n4474,n4473);
and gate_3974(n4475,n4466,n4474);
not gate_3975(po112,n4475);
and gate_3976(n4477,pi131,n629);
not gate_3977(n4478,n4477);
and gate_3978(n4479,pi116,pi198);
not gate_3979(n4480,n4479);
and gate_3980(n4481,pi124,n570);
not gate_3981(n4482,n4481);
and gate_3982(n4483,n4480,n4482);
not gate_3983(n4484,n4483);
and gate_3984(n4485,n630,n4484);
not gate_3985(n4486,n4485);
and gate_3986(n4487,n4478,n4486);
not gate_3987(po113,n4487);
and gate_3988(n4489,n3662,n4038);
and gate_3989(n4490,n3658,n4489);
and gate_3990(n4491,n3673,n4035);
and gate_3991(n4492,n3621,n4024);
not gate_3992(n4493,n4492);
and gate_3993(n4494,n3688,n4493);
and gate_3994(n4495,n4491,n4494);
and gate_3995(n4496,n4490,n4495);
and gate_3996(n4497,n3694,n4021);
and gate_3997(n4498,n4019,n4497);
and gate_3998(n4499,n3622,n3686);
not gate_3999(n4500,n4499);
and gate_4000(n4501,n3696,n4500);
and gate_4001(n4502,n3706,n4501);
and gate_4002(n4503,n4498,n4502);
and gate_4003(n4504,n4496,n4503);
and gate_4004(n4505,n3621,n3770);
not gate_4005(n4506,n4505);
and gate_4006(n4507,n3736,n4506);
and gate_4007(n4508,n3730,n4507);
and gate_4008(n4509,n4048,n4508);
and gate_4009(n4510,n3757,n4065);
and gate_4010(n4511,n4063,n4510);
and gate_4011(n4512,n3768,n3775);
and gate_4012(n4513,n3622,n3732);
not gate_4013(n4514,n4513);
and gate_4014(n4515,n3795,n4033);
not gate_4015(n4516,n4515);
and gate_4016(n4517,n4514,n4516);
and gate_4017(n4518,n4512,n4517);
and gate_4018(n4519,n4511,n4518);
and gate_4019(n4520,n4509,n4519);
and gate_4020(n4521,n4504,n4520);
and gate_4021(n4522,n3634,n3674);
and gate_4022(n4523,n3678,n4522);
not gate_4023(n4524,n4523);
and gate_4024(n4525,n3621,n3634);
not gate_4025(n4526,n4525);
and gate_4026(n4527,n3796,n4526);
not gate_4027(n4528,n4527);
and gate_4028(n4529,n3627,n4527);
and gate_4029(n4530,n3739,n4529);
not gate_4030(n4531,n4530);
and gate_4031(n4532,n4524,n4531);
not gate_4032(n4533,n4532);
and gate_4033(n4534,n3640,n4533);
not gate_4034(n4535,n4534);
and gate_4035(n4536,n4521,n4535);
not gate_4036(n4537,n4536);
and gate_4037(n4538,n543,n4537);
not gate_4038(n4539,n4538);
and gate_4039(n4540,pi171,n4536);
not gate_4040(n4541,n4540);
and gate_4041(n4542,n4539,n4541);
not gate_4042(n4543,n4542);
and gate_4043(n4544,n629,n4543);
not gate_4044(n4545,n4544);
and gate_4045(n4546,pi117,pi198);
not gate_4046(n4547,n4546);
and gate_4047(n4548,pi125,n570);
not gate_4048(n4549,n4548);
and gate_4049(n4550,n4547,n4549);
not gate_4050(n4551,n4550);
and gate_4051(n4552,n630,n4551);
not gate_4052(n4553,n4552);
and gate_4053(n4554,n4545,n4553);
not gate_4054(po114,n4554);
and gate_4055(n4556,pi139,n629);
not gate_4056(n4557,n4556);
and gate_4057(n4558,pi118,pi198);
not gate_4058(n4559,n4558);
and gate_4059(n4560,pi126,n570);
not gate_4060(n4561,n4560);
and gate_4061(n4562,n4559,n4561);
not gate_4062(n4563,n4562);
and gate_4063(n4564,n630,n4563);
not gate_4064(n4565,n4564);
and gate_4065(n4566,n4557,n4565);
not gate_4066(po115,n4566);
and gate_4067(n4568,n4075,n4528);
and gate_4068(n4569,n3627,n4568);
and gate_4069(n4570,n3639,n4569);
and gate_4070(n4571,n3646,n4570);
not gate_4071(n4572,n4571);
and gate_4072(n4573,n3683,n4493);
and gate_4073(n4574,n4036,n4573);
and gate_4074(n4575,n3668,n3673);
and gate_4075(n4576,n4574,n4575);
and gate_4076(n4577,n3714,n4019);
and gate_4077(n4578,n3705,n4026);
and gate_4078(n4579,n4501,n4578);
and gate_4079(n4580,n4577,n4579);
and gate_4080(n4581,n4576,n4580);
and gate_4081(n4582,n3750,n4047);
and gate_4082(n4583,n4052,n4507);
and gate_4083(n4584,n4582,n4583);
and gate_4084(n4585,n3762,n4065);
and gate_4085(n4586,n4056,n4514);
and gate_4086(n4587,n3769,n4586);
and gate_4087(n4588,n4585,n4587);
and gate_4088(n4589,n4584,n4588);
and gate_4089(n4590,n4581,n4589);
and gate_4090(n4591,n3628,n4076);
and gate_4091(n4592,n3633,n4591);
and gate_4092(n4593,n3640,n4592);
and gate_4093(n4594,n3645,n4593);
not gate_4094(n4595,n4594);
and gate_4095(n4596,n4590,n4595);
and gate_4096(n4597,n4572,n4596);
not gate_4097(n4598,n4597);
and gate_4098(n4599,n551,n4598);
not gate_4099(n4600,n4599);
and gate_4100(n4601,pi179,n4597);
not gate_4101(n4602,n4601);
and gate_4102(n4603,n4600,n4602);
not gate_4103(n4604,n4603);
and gate_4104(n4605,n629,n4604);
not gate_4105(n4606,n4605);
and gate_4106(n4607,pi119,pi198);
not gate_4107(n4608,n4607);
and gate_4108(n4609,pi127,n570);
not gate_4109(n4610,n4609);
and gate_4110(n4611,n4608,n4610);
not gate_4111(n4612,n4611);
and gate_4112(n4613,n630,n4612);
not gate_4113(n4614,n4613);
and gate_4114(n4615,n4606,n4614);
not gate_4115(po116,n4615);
and gate_4116(n4617,pi147,n629);
not gate_4117(n4618,n4617);
and gate_4118(n4619,pi120,pi198);
not gate_4119(n4620,n4619);
and gate_4120(n4621,pi128,n570);
not gate_4121(n4622,n4621);
and gate_4122(n4623,n4620,n4622);
not gate_4123(n4624,n4623);
and gate_4124(n4625,n630,n4624);
not gate_4125(n4626,n4625);
and gate_4126(n4627,n4618,n4626);
not gate_4127(po117,n4627);
and gate_4128(n4629,n1063,n3935);
and gate_4129(n4630,n1075,n2780);
and gate_4130(n4631,n3940,n4630);
and gate_4131(n4632,n4629,n4631);
and gate_4132(n4633,n1088,n3946);
and gate_4133(n4634,n1094,n4633);
and gate_4134(n4635,n1098,n2793);
and gate_4135(n4636,n1105,n2789);
and gate_4136(n4637,n4635,n4636);
and gate_4137(n4638,n4634,n4637);
and gate_4138(n4639,n4632,n4638);
and gate_4139(n4640,n1123,n2798);
and gate_4140(n4641,n1119,n4640);
and gate_4141(n4642,n1138,n3954);
and gate_4142(n4643,n2807,n4642);
and gate_4143(n4644,n4641,n4643);
and gate_4144(n4645,n1159,n3966);
and gate_4145(n4646,n1162,n2811);
and gate_4146(n4647,n2819,n4646);
and gate_4147(n4648,n4645,n4647);
and gate_4148(n4649,n4644,n4648);
and gate_4149(n4650,n4639,n4649);
and gate_4150(n4651,n1188,n2759);
and gate_4151(n4652,n1071,n4651);
not gate_4152(n4653,n4652);
and gate_4153(n4654,n4650,n4653);
and gate_4154(n4655,n1028,n1176);
and gate_4155(n4656,n1034,n1039);
not gate_4156(n4657,n4656);
and gate_4157(n4658,n2755,n4657);
and gate_4158(n4659,n4655,n4658);
and gate_4159(n4660,n1114,n4659);
not gate_4160(n4661,n4660);
and gate_4161(n4662,n4654,n4661);
not gate_4162(n4663,n4662);
and gate_4163(n4664,n559,n4663);
not gate_4164(n4665,n4664);
and gate_4165(n4666,pi187,n4662);
not gate_4166(n4667,n4666);
and gate_4167(n4668,n4665,n4667);
not gate_4168(n4669,n4668);
and gate_4169(n4670,n629,n4669);
not gate_4170(n4671,n4670);
and gate_4171(n4672,pi129,n570);
not gate_4172(n4673,n4672);
and gate_4173(n4674,pi121,pi198);
not gate_4174(n4675,n4674);
and gate_4175(n4676,n4673,n4675);
not gate_4176(n4677,n4676);
and gate_4177(n4678,n630,n4677);
not gate_4178(n4679,n4678);
and gate_4179(n4680,n4671,n4679);
not gate_4180(po118,n4680);
and gate_4181(n4682,pi155,n629);
not gate_4182(n4683,n4682);
and gate_4183(n4684,pi130,n570);
not gate_4184(n4685,n4684);
and gate_4185(n4686,pi122,pi198);
not gate_4186(n4687,n4686);
and gate_4187(n4688,n4685,n4687);
not gate_4188(n4689,n4688);
and gate_4189(n4690,n630,n4689);
not gate_4190(n4691,n4690);
and gate_4191(n4692,n4683,n4691);
not gate_4192(po119,n4692);
and gate_4193(n4694,n630,n4464);
not gate_4194(n4695,n4694);
and gate_4195(n4696,pi001,n629);
not gate_4196(n4697,n4696);
and gate_4197(n4698,n4695,n4697);
not gate_4198(po120,n4698);
and gate_4199(n4700,n630,n4176);
not gate_4200(n4701,n4700);
and gate_4201(n4702,pi060,n629);
not gate_4202(n4703,n4702);
and gate_4203(n4704,n4701,n4703);
not gate_4204(po121,n4704);
and gate_4205(n4706,n630,n3811);
not gate_4206(n4707,n4706);
and gate_4207(n4708,pi052,n629);
not gate_4208(n4709,n4708);
and gate_4209(n4710,n4707,n4709);
not gate_4210(po122,n4710);
and gate_4211(n4712,n630,n3333);
not gate_4212(n4713,n4712);
and gate_4213(n4714,pi044,n629);
not gate_4214(n4715,n4714);
and gate_4215(n4716,n4713,n4715);
not gate_4216(po123,n4716);
and gate_4217(n4718,n630,n2902);
not gate_4218(n4719,n4718);
and gate_4219(n4720,pi036,n629);
not gate_4220(n4721,n4720);
and gate_4221(n4722,n4719,n4721);
not gate_4222(po124,n4722);
and gate_4223(n4724,n630,n2420);
not gate_4224(n4725,n4724);
and gate_4225(n4726,pi028,n629);
not gate_4226(n4727,n4726);
and gate_4227(n4728,n4725,n4727);
not gate_4228(po125,n4728);
and gate_4229(n4730,n630,n1799);
not gate_4230(n4731,n4730);
and gate_4231(n4732,pi020,n629);
not gate_4232(n4733,n4732);
and gate_4233(n4734,n4731,n4733);
not gate_4234(po126,n4734);
and gate_4235(n4736,n630,n1203);
not gate_4236(n4737,n4736);
and gate_4237(n4738,pi012,n629);
not gate_4238(n4739,n4738);
and gate_4239(n4740,n4737,n4739);
not gate_4240(po127,n4740);
and gate_4241(n4742,n630,n4543);
not gate_4242(n4743,n4742);
and gate_4243(n4744,pi003,n629);
not gate_4244(n4745,n4744);
and gate_4245(n4746,n4743,n4745);
not gate_4246(po128,n4746);
and gate_4247(n4748,n630,n4240);
not gate_4248(n4749,n4748);
and gate_4249(n4750,pi062,n629);
not gate_4250(n4751,n4750);
and gate_4251(n4752,n4749,n4751);
not gate_4252(po129,n4752);
and gate_4253(n4754,n630,n3909);
not gate_4254(n4755,n4754);
and gate_4255(n4756,pi054,n629);
not gate_4256(n4757,n4756);
and gate_4257(n4758,n4755,n4757);
not gate_4258(po130,n4758);
and gate_4259(n4760,n630,n3434);
not gate_4260(n4761,n4760);
and gate_4261(n4762,pi046,n629);
not gate_4262(n4763,n4762);
and gate_4263(n4764,n4761,n4763);
not gate_4264(po131,n4764);
and gate_4265(n4766,n630,n2967);
not gate_4266(n4767,n4766);
and gate_4267(n4768,pi038,n629);
not gate_4268(n4769,n4768);
and gate_4269(n4770,n4767,n4769);
not gate_4270(po132,n4770);
and gate_4271(n4772,n630,n2637);
not gate_4272(n4773,n4772);
and gate_4273(n4774,pi030,n629);
not gate_4274(n4775,n4774);
and gate_4275(n4776,n4773,n4775);
not gate_4276(po133,n4776);
and gate_4277(n4778,n630,n2023);
not gate_4278(n4779,n4778);
and gate_4279(n4780,pi022,n629);
not gate_4280(n4781,n4780);
and gate_4281(n4782,n4779,n4781);
not gate_4282(po134,n4782);
and gate_4283(n4784,n630,n1412);
not gate_4284(n4785,n4784);
and gate_4285(n4786,pi014,n629);
not gate_4286(n4787,n4786);
and gate_4287(n4788,n4785,n4787);
not gate_4288(po135,n4788);
and gate_4289(n4790,n630,n4604);
not gate_4290(n4791,n4790);
and gate_4291(n4792,pi005,n629);
not gate_4292(n4793,n4792);
and gate_4293(n4794,n4791,n4793);
not gate_4294(po136,n4794);
and gate_4295(n4796,n630,n4313);
not gate_4296(n4797,n4796);
and gate_4297(n4798,pi064,n629);
not gate_4298(n4799,n4798);
and gate_4299(n4800,n4797,n4799);
not gate_4300(po137,n4800);
and gate_4301(n4802,n630,n3993);
not gate_4302(n4803,n4802);
and gate_4303(n4804,pi056,n629);
not gate_4304(n4805,n4804);
and gate_4305(n4806,n4803,n4805);
not gate_4306(po138,n4806);
and gate_4307(n4808,n630,n3516);
not gate_4308(n4809,n4808);
and gate_4309(n4810,pi048,n629);
not gate_4310(n4811,n4810);
and gate_4311(n4812,n4809,n4811);
not gate_4312(po139,n4812);
and gate_4313(n4814,n630,n3179);
not gate_4314(n4815,n4814);
and gate_4315(n4816,pi040,n629);
not gate_4316(n4817,n4816);
and gate_4317(n4818,n4815,n4817);
not gate_4318(po140,n4818);
and gate_4319(n4820,n630,n2729);
not gate_4320(n4821,n4820);
and gate_4321(n4822,pi032,n629);
not gate_4322(n4823,n4822);
and gate_4323(n4824,n4821,n4823);
not gate_4324(po141,n4824);
and gate_4325(n4826,n630,n2101);
not gate_4326(n4827,n4826);
and gate_4327(n4828,pi024,n629);
not gate_4328(n4829,n4828);
and gate_4329(n4830,n4827,n4829);
not gate_4330(po142,n4830);
and gate_4331(n4832,n630,n1502);
not gate_4332(n4833,n4832);
and gate_4333(n4834,pi016,n629);
not gate_4334(n4835,n4834);
and gate_4335(n4836,n4833,n4835);
not gate_4336(po143,n4836);
and gate_4337(n4838,n630,n4669);
not gate_4338(n4839,n4838);
and gate_4339(n4840,pi007,n629);
not gate_4340(n4841,n4840);
and gate_4341(n4842,n4839,n4841);
not gate_4342(po144,n4842);
and gate_4343(n4844,n630,n4393);
not gate_4344(n4845,n4844);
and gate_4345(n4846,pi066,n629);
not gate_4346(n4847,n4846);
and gate_4347(n4848,n4845,n4847);
not gate_4348(po145,n4848);
and gate_4349(n4850,n630,n4095);
not gate_4350(n4851,n4850);
and gate_4351(n4852,pi058,n629);
not gate_4352(n4853,n4852);
and gate_4353(n4854,n4851,n4853);
not gate_4354(po146,n4854);
and gate_4355(n4856,n630,n3592);
not gate_4356(n4857,n4856);
and gate_4357(n4858,pi050,n629);
not gate_4358(n4859,n4858);
and gate_4359(n4860,n4857,n4859);
not gate_4360(po147,n4860);
and gate_4361(n4862,n630,n3266);
not gate_4362(n4863,n4862);
and gate_4363(n4864,pi042,n629);
not gate_4364(n4865,n4864);
and gate_4365(n4866,n4863,n4865);
not gate_4366(po148,n4866);
and gate_4367(n4868,n630,n2834);
not gate_4368(n4869,n4868);
and gate_4369(n4870,pi034,n629);
not gate_4370(n4871,n4870);
and gate_4371(n4872,n4869,n4871);
not gate_4372(po149,n4872);
and gate_4373(n4874,n630,n2200);
not gate_4374(n4875,n4874);
and gate_4375(n4876,pi026,n629);
not gate_4376(n4877,n4876);
and gate_4377(n4878,n4875,n4877);
not gate_4378(po150,n4878);
and gate_4379(n4880,n630,n1708);
not gate_4380(n4881,n4880);
and gate_4381(n4882,pi018,n629);
not gate_4382(n4883,n4882);
and gate_4383(n4884,n4881,n4883);
not gate_4384(po151,n4884);
and gate_4385(n4886,pi131,n630);
not gate_4386(n4887,n4886);
and gate_4387(n4888,pi000,n629);
not gate_4388(n4889,n4888);
and gate_4389(n4890,n4887,n4889);
not gate_4390(po152,n4890);
and gate_4391(n4892,pi132,n630);
not gate_4392(n4893,n4892);
and gate_4393(n4894,pi059,n629);
not gate_4394(n4895,n4894);
and gate_4395(n4896,n4893,n4895);
not gate_4396(po153,n4896);
and gate_4397(n4898,pi133,n630);
not gate_4398(n4899,n4898);
and gate_4399(n4900,pi051,n629);
not gate_4400(n4901,n4900);
and gate_4401(n4902,n4899,n4901);
not gate_4402(po154,n4902);
and gate_4403(n4904,pi134,n630);
not gate_4404(n4905,n4904);
and gate_4405(n4906,pi043,n629);
not gate_4406(n4907,n4906);
and gate_4407(n4908,n4905,n4907);
not gate_4408(po155,n4908);
and gate_4409(n4910,pi135,n630);
not gate_4410(n4911,n4910);
and gate_4411(n4912,pi035,n629);
not gate_4412(n4913,n4912);
and gate_4413(n4914,n4911,n4913);
not gate_4414(po156,n4914);
and gate_4415(n4916,pi136,n630);
not gate_4416(n4917,n4916);
and gate_4417(n4918,pi027,n629);
not gate_4418(n4919,n4918);
and gate_4419(n4920,n4917,n4919);
not gate_4420(po157,n4920);
and gate_4421(n4922,pi137,n630);
not gate_4422(n4923,n4922);
and gate_4423(n4924,pi019,n629);
not gate_4424(n4925,n4924);
and gate_4425(n4926,n4923,n4925);
not gate_4426(po158,n4926);
and gate_4427(n4928,pi138,n630);
not gate_4428(n4929,n4928);
and gate_4429(n4930,pi011,n629);
not gate_4430(n4931,n4930);
and gate_4431(n4932,n4929,n4931);
not gate_4432(po159,n4932);
and gate_4433(n4934,pi139,n630);
not gate_4434(n4935,n4934);
and gate_4435(n4936,pi002,n629);
not gate_4436(n4937,n4936);
and gate_4437(n4938,n4935,n4937);
not gate_4438(po160,n4938);
and gate_4439(n4940,pi140,n630);
not gate_4440(n4941,n4940);
and gate_4441(n4942,pi061,n629);
not gate_4442(n4943,n4942);
and gate_4443(n4944,n4941,n4943);
not gate_4444(po161,n4944);
and gate_4445(n4946,pi141,n630);
not gate_4446(n4947,n4946);
and gate_4447(n4948,pi053,n629);
not gate_4448(n4949,n4948);
and gate_4449(n4950,n4947,n4949);
not gate_4450(po162,n4950);
and gate_4451(n4952,pi142,n630);
not gate_4452(n4953,n4952);
and gate_4453(n4954,pi045,n629);
not gate_4454(n4955,n4954);
and gate_4455(n4956,n4953,n4955);
not gate_4456(po163,n4956);
and gate_4457(n4958,pi143,n630);
not gate_4458(n4959,n4958);
and gate_4459(n4960,pi037,n629);
not gate_4460(n4961,n4960);
and gate_4461(n4962,n4959,n4961);
not gate_4462(po164,n4962);
and gate_4463(n4964,pi144,n630);
not gate_4464(n4965,n4964);
and gate_4465(n4966,pi029,n629);
not gate_4466(n4967,n4966);
and gate_4467(n4968,n4965,n4967);
not gate_4468(po165,n4968);
and gate_4469(n4970,pi145,n630);
not gate_4470(n4971,n4970);
and gate_4471(n4972,pi021,n629);
not gate_4472(n4973,n4972);
and gate_4473(n4974,n4971,n4973);
not gate_4474(po166,n4974);
and gate_4475(n4976,pi146,n630);
not gate_4476(n4977,n4976);
and gate_4477(n4978,pi013,n629);
not gate_4478(n4979,n4978);
and gate_4479(n4980,n4977,n4979);
not gate_4480(po167,n4980);
and gate_4481(n4982,pi147,n630);
not gate_4482(n4983,n4982);
and gate_4483(n4984,pi004,n629);
not gate_4484(n4985,n4984);
and gate_4485(n4986,n4983,n4985);
not gate_4486(po168,n4986);
and gate_4487(n4988,pi148,n630);
not gate_4488(n4989,n4988);
and gate_4489(n4990,pi063,n629);
not gate_4490(n4991,n4990);
and gate_4491(n4992,n4989,n4991);
not gate_4492(po169,n4992);
and gate_4493(n4994,pi149,n630);
not gate_4494(n4995,n4994);
and gate_4495(n4996,pi055,n629);
not gate_4496(n4997,n4996);
and gate_4497(n4998,n4995,n4997);
not gate_4498(po170,n4998);
and gate_4499(n5000,pi150,n630);
not gate_4500(n5001,n5000);
and gate_4501(n5002,pi047,n629);
not gate_4502(n5003,n5002);
and gate_4503(n5004,n5001,n5003);
not gate_4504(po171,n5004);
and gate_4505(n5006,pi151,n630);
not gate_4506(n5007,n5006);
and gate_4507(n5008,pi039,n629);
not gate_4508(n5009,n5008);
and gate_4509(n5010,n5007,n5009);
not gate_4510(po172,n5010);
and gate_4511(n5012,pi152,n630);
not gate_4512(n5013,n5012);
and gate_4513(n5014,pi031,n629);
not gate_4514(n5015,n5014);
and gate_4515(n5016,n5013,n5015);
not gate_4516(po173,n5016);
and gate_4517(n5018,pi153,n630);
not gate_4518(n5019,n5018);
and gate_4519(n5020,pi023,n629);
not gate_4520(n5021,n5020);
and gate_4521(n5022,n5019,n5021);
not gate_4522(po174,n5022);
and gate_4523(n5024,pi154,n630);
not gate_4524(n5025,n5024);
and gate_4525(n5026,pi015,n629);
not gate_4526(n5027,n5026);
and gate_4527(n5028,n5025,n5027);
not gate_4528(po175,n5028);
and gate_4529(n5030,pi155,n630);
not gate_4530(n5031,n5030);
and gate_4531(n5032,pi006,n629);
not gate_4532(n5033,n5032);
and gate_4533(n5034,n5031,n5033);
not gate_4534(po176,n5034);
and gate_4535(n5036,pi156,n630);
not gate_4536(n5037,n5036);
and gate_4537(n5038,pi065,n629);
not gate_4538(n5039,n5038);
and gate_4539(n5040,n5037,n5039);
not gate_4540(po177,n5040);
and gate_4541(n5042,pi157,n630);
not gate_4542(n5043,n5042);
and gate_4543(n5044,pi057,n629);
not gate_4544(n5045,n5044);
and gate_4545(n5046,n5043,n5045);
not gate_4546(po178,n5046);
and gate_4547(n5048,pi158,n630);
not gate_4548(n5049,n5048);
and gate_4549(n5050,pi049,n629);
not gate_4550(n5051,n5050);
and gate_4551(n5052,n5049,n5051);
not gate_4552(po179,n5052);
and gate_4553(n5054,pi159,n630);
not gate_4554(n5055,n5054);
and gate_4555(n5056,pi041,n629);
not gate_4556(n5057,n5056);
and gate_4557(n5058,n5055,n5057);
not gate_4558(po180,n5058);
and gate_4559(n5060,pi160,n630);
not gate_4560(n5061,n5060);
and gate_4561(n5062,pi033,n629);
not gate_4562(n5063,n5062);
and gate_4563(n5064,n5061,n5063);
not gate_4564(po181,n5064);
and gate_4565(n5066,pi161,n630);
not gate_4566(n5067,n5066);
and gate_4567(n5068,pi025,n629);
not gate_4568(n5069,n5068);
and gate_4569(n5070,n5067,n5069);
not gate_4570(po182,n5070);
and gate_4571(n5072,pi162,n630);
not gate_4572(n5073,n5072);
and gate_4573(n5074,pi017,n629);
not gate_4574(n5075,n5074);
and gate_4575(n5076,n5073,n5075);
not gate_4576(po183,n5076);
and gate_4577(n5078,pi196,n626);
not gate_4578(n5079,n5078);
and gate_4579(n5080,pi195,n5079);
not gate_4580(n5081,n5080);
and gate_4581(n5082,n567,n5078);
not gate_4582(n5083,n5082);
and gate_4583(n5084,n5081,n5083);
not gate_4584(n5085,n5084);
and gate_4585(n5086,pi010,n629);
not gate_4586(n5087,n5086);
and gate_4587(n5088,n501,n5087);
and gate_4588(po184,n5085,n5088);
and gate_4589(n5090,n568,n627);
not gate_4590(n5091,n5090);
and gate_4591(n5092,n5079,n5091);
and gate_4592(po185,n5088,n5092);
and gate_4593(n5094,pi197,n570);
not gate_4594(n5095,n5094);
and gate_4595(n5096,n569,pi198);
not gate_4596(n5097,n5096);
and gate_4597(n5098,n5095,n5097);
not gate_4598(n5099,n5098);
and gate_4599(po186,n5088,n5099);
and gate_4600(po187,n570,n5088);
and gate_4601(n5102,n502,pi039);
not gate_4602(n5103,n5102);
and gate_4603(n5104,pi009,pi018);
not gate_4604(n5105,n5104);
and gate_4605(n5106,n5103,n5105);
not gate_4606(n5107,n5106);
and gate_4607(n5108,n5086,n5107);
not gate_4608(n5109,n5108);
and gate_4609(n5110,pi196,pi197);
and gate_4610(n5111,n567,n570);
not gate_4611(n5112,n5111);
and gate_4612(n5113,n5110,n5112);
not gate_4613(n5114,n5113);
and gate_4614(n5115,n568,n569);
and gate_4615(n5116,n5111,n5115);
not gate_4616(n5117,n5116);
and gate_4617(n5118,n5114,n5117);
not gate_4618(n5119,n5118);
and gate_4619(n5120,pi226,n5119);
not gate_4620(n5121,n5120);
and gate_4621(n5122,pi225,n5118);
not gate_4622(n5123,n5122);
and gate_4623(n5124,n5121,n5123);
not gate_4624(n5125,n5124);
and gate_4625(n5126,pi255,n5125);
not gate_4626(n5127,n5126);
and gate_4627(n5128,pi200,n5119);
not gate_4628(n5129,n5128);
and gate_4629(n5130,pi201,n5118);
not gate_4630(n5131,n5130);
and gate_4631(n5132,n5129,n5131);
not gate_4632(n5133,n5132);
and gate_4633(n5134,n619,n5133);
not gate_4634(n5135,n5134);
and gate_4635(n5136,n5127,n5135);
not gate_4636(n5137,n5136);
and gate_4637(n5138,n502,pi255);
not gate_4638(n5139,n5138);
and gate_4639(n5140,pi009,n619);
not gate_4640(n5141,n5140);
and gate_4641(n5142,n5139,n5141);
not gate_4642(n5143,n5142);
and gate_4643(n5144,n629,n5143);
not gate_4644(n5145,n5144);
and gate_4645(n5146,n5137,n5145);
not gate_4646(n5147,n5146);
and gate_4647(n5148,pi199,n5144);
not gate_4648(n5149,n5148);
and gate_4649(n5150,n5147,n5149);
not gate_4650(n5151,n5150);
and gate_4651(n5152,n5087,n5151);
not gate_4652(n5153,n5152);
and gate_4653(n5154,n5109,n5153);
not gate_4654(n5155,n5154);
and gate_4655(po188,n501,n5155);
and gate_4656(n5157,pi009,pi039);
not gate_4657(n5158,n5157);
and gate_4658(n5159,n502,pi031);
not gate_4659(n5160,n5159);
and gate_4660(n5161,n5158,n5160);
not gate_4661(n5162,n5161);
and gate_4662(n5163,n5086,n5162);
not gate_4663(n5164,n5163);
and gate_4664(n5165,pi199,n5119);
not gate_4665(n5166,n5165);
and gate_4666(n5167,pi226,n5118);
not gate_4667(n5168,n5167);
and gate_4668(n5169,n5166,n5168);
not gate_4669(n5170,n5169);
and gate_4670(n5171,pi255,n5170);
not gate_4671(n5172,n5171);
and gate_4672(n5173,pi201,n5119);
not gate_4673(n5174,n5173);
and gate_4674(n5175,pi202,n5118);
not gate_4675(n5176,n5175);
and gate_4676(n5177,n5174,n5176);
not gate_4677(n5178,n5177);
and gate_4678(n5179,n619,n5178);
not gate_4679(n5180,n5179);
and gate_4680(n5181,n5172,n5180);
not gate_4681(n5182,n5181);
and gate_4682(n5183,n5145,n5182);
not gate_4683(n5184,n5183);
and gate_4684(n5185,pi200,n5144);
not gate_4685(n5186,n5185);
and gate_4686(n5187,n5184,n5186);
not gate_4687(n5188,n5187);
and gate_4688(n5189,n5087,n5188);
not gate_4689(n5190,n5189);
and gate_4690(n5191,n5164,n5190);
not gate_4691(n5192,n5191);
and gate_4692(po189,n501,n5192);
and gate_4693(n5194,pi199,n5118);
not gate_4694(n5195,n5194);
and gate_4695(n5196,n5129,n5195);
not gate_4696(n5197,n5196);
and gate_4697(n5198,pi255,n5197);
not gate_4698(n5199,n5198);
and gate_4699(n5200,pi202,n5119);
not gate_4700(n5201,n5200);
and gate_4701(n5202,pi203,n5118);
not gate_4702(n5203,n5202);
and gate_4703(n5204,n5201,n5203);
not gate_4704(n5205,n5204);
and gate_4705(n5206,n619,n5205);
not gate_4706(n5207,n5206);
and gate_4707(n5208,n5199,n5207);
not gate_4708(n5209,n5208);
and gate_4709(n5210,n5145,n5209);
not gate_4710(n5211,n5210);
and gate_4711(n5212,pi201,n5144);
not gate_4712(n5213,n5212);
and gate_4713(n5214,n5211,n5213);
not gate_4714(n5215,n5214);
and gate_4715(n5216,n5087,n5215);
not gate_4716(n5217,n5216);
and gate_4717(n5218,pi009,pi031);
not gate_4718(n5219,n5218);
and gate_4719(n5220,n502,pi023);
not gate_4720(n5221,n5220);
and gate_4721(n5222,n5219,n5221);
not gate_4722(n5223,n5222);
and gate_4723(n5224,n5086,n5223);
not gate_4724(n5225,n5224);
and gate_4725(n5226,n5217,n5225);
not gate_4726(n5227,n5226);
and gate_4727(po190,n501,n5227);
and gate_4728(n5229,pi200,n5118);
not gate_4729(n5230,n5229);
and gate_4730(n5231,n5174,n5230);
not gate_4731(n5232,n5231);
and gate_4732(n5233,pi255,n5232);
not gate_4733(n5234,n5233);
and gate_4734(n5235,pi203,n5119);
not gate_4735(n5236,n5235);
and gate_4736(n5237,pi204,n5118);
not gate_4737(n5238,n5237);
and gate_4738(n5239,n5236,n5238);
not gate_4739(n5240,n5239);
and gate_4740(n5241,n619,n5240);
not gate_4741(n5242,n5241);
and gate_4742(n5243,n5234,n5242);
not gate_4743(n5244,n5243);
and gate_4744(n5245,n5145,n5244);
not gate_4745(n5246,n5245);
and gate_4746(n5247,pi202,n5144);
not gate_4747(n5248,n5247);
and gate_4748(n5249,n5246,n5248);
not gate_4749(n5250,n5249);
and gate_4750(n5251,n5087,n5250);
not gate_4751(n5252,n5251);
and gate_4752(n5253,pi009,pi023);
not gate_4753(n5254,n5253);
and gate_4754(n5255,n502,pi015);
not gate_4755(n5256,n5255);
and gate_4756(n5257,n5254,n5256);
not gate_4757(n5258,n5257);
and gate_4758(n5259,n5086,n5258);
not gate_4759(n5260,n5259);
and gate_4760(n5261,n5252,n5260);
not gate_4761(n5262,n5261);
and gate_4762(po191,n501,n5262);
and gate_4763(n5264,pi005,n502);
not gate_4764(n5265,n5264);
and gate_4765(n5266,pi009,pi015);
not gate_4766(n5267,n5266);
and gate_4767(n5268,n5265,n5267);
not gate_4768(n5269,n5268);
and gate_4769(n5270,n5086,n5269);
not gate_4770(n5271,n5270);
and gate_4771(n5272,n5131,n5201);
not gate_4772(n5273,n5272);
and gate_4773(n5274,pi255,n5273);
not gate_4774(n5275,n5274);
and gate_4775(n5276,pi205,n5118);
not gate_4776(n5277,n5276);
and gate_4777(n5278,pi204,n5119);
not gate_4778(n5279,n5278);
and gate_4779(n5280,n5277,n5279);
not gate_4780(n5281,n5280);
and gate_4781(n5282,n619,n5281);
not gate_4782(n5283,n5282);
and gate_4783(n5284,n5275,n5283);
not gate_4784(n5285,n5284);
and gate_4785(n5286,n5145,n5285);
not gate_4786(n5287,n5286);
and gate_4787(n5288,pi203,n5144);
not gate_4788(n5289,n5288);
and gate_4789(n5290,n5287,n5289);
not gate_4790(n5291,n5290);
and gate_4791(n5292,n5087,n5291);
not gate_4792(n5293,n5292);
and gate_4793(n5294,n5271,n5293);
not gate_4794(n5295,n5294);
and gate_4795(po192,n501,n5295);
and gate_4796(n5297,pi005,pi009);
not gate_4797(n5298,n5297);
and gate_4798(n5299,n502,pi064);
not gate_4799(n5300,n5299);
and gate_4800(n5301,n5298,n5300);
not gate_4801(n5302,n5301);
and gate_4802(n5303,n5086,n5302);
not gate_4803(n5304,n5303);
and gate_4804(n5305,n5176,n5236);
not gate_4805(n5306,n5305);
and gate_4806(n5307,pi255,n5306);
not gate_4807(n5308,n5307);
and gate_4808(n5309,pi206,n5118);
not gate_4809(n5310,n5309);
and gate_4810(n5311,pi205,n5119);
not gate_4811(n5312,n5311);
and gate_4812(n5313,n5310,n5312);
not gate_4813(n5314,n5313);
and gate_4814(n5315,n619,n5314);
not gate_4815(n5316,n5315);
and gate_4816(n5317,n5308,n5316);
not gate_4817(n5318,n5317);
and gate_4818(n5319,n5145,n5318);
not gate_4819(n5320,n5319);
and gate_4820(n5321,pi204,n5144);
not gate_4821(n5322,n5321);
and gate_4822(n5323,n5320,n5322);
not gate_4823(n5324,n5323);
and gate_4824(n5325,n5087,n5324);
not gate_4825(n5326,n5325);
and gate_4826(n5327,n5304,n5326);
not gate_4827(n5328,n5327);
and gate_4828(po193,n501,n5328);
and gate_4829(n5330,n502,pi056);
not gate_4830(n5331,n5330);
and gate_4831(n5332,pi009,pi064);
not gate_4832(n5333,n5332);
and gate_4833(n5334,n5331,n5333);
not gate_4834(n5335,n5334);
and gate_4835(n5336,n5086,n5335);
not gate_4836(n5337,n5336);
and gate_4837(n5338,n5203,n5279);
not gate_4838(n5339,n5338);
and gate_4839(n5340,pi255,n5339);
not gate_4840(n5341,n5340);
and gate_4841(n5342,pi206,n5119);
not gate_4842(n5343,n5342);
and gate_4843(n5344,pi207,n5118);
not gate_4844(n5345,n5344);
and gate_4845(n5346,n5343,n5345);
not gate_4846(n5347,n5346);
and gate_4847(n5348,n619,n5347);
not gate_4848(n5349,n5348);
and gate_4849(n5350,n5341,n5349);
not gate_4850(n5351,n5350);
and gate_4851(n5352,n5145,n5351);
not gate_4852(n5353,n5352);
and gate_4853(n5354,pi205,n5144);
not gate_4854(n5355,n5354);
and gate_4855(n5356,n5353,n5355);
not gate_4856(n5357,n5356);
and gate_4857(n5358,n5087,n5357);
not gate_4858(n5359,n5358);
and gate_4859(n5360,n5337,n5359);
not gate_4860(n5361,n5360);
and gate_4861(po194,n501,n5361);
and gate_4862(n5363,n5238,n5312);
not gate_4863(n5364,n5363);
and gate_4864(n5365,pi255,n5364);
not gate_4865(n5366,n5365);
and gate_4866(n5367,pi207,n5119);
not gate_4867(n5368,n5367);
and gate_4868(n5369,pi208,n5118);
not gate_4869(n5370,n5369);
and gate_4870(n5371,n5368,n5370);
not gate_4871(n5372,n5371);
and gate_4872(n5373,n619,n5372);
not gate_4873(n5374,n5373);
and gate_4874(n5375,n5366,n5374);
not gate_4875(n5376,n5375);
and gate_4876(n5377,n5145,n5376);
not gate_4877(n5378,n5377);
and gate_4878(n5379,pi206,n5144);
not gate_4879(n5380,n5379);
and gate_4880(n5381,n5378,n5380);
not gate_4881(n5382,n5381);
and gate_4882(n5383,n5087,n5382);
not gate_4883(n5384,n5383);
and gate_4884(n5385,pi009,pi056);
not gate_4885(n5386,n5385);
and gate_4886(n5387,n502,pi048);
not gate_4887(n5388,n5387);
and gate_4888(n5389,n5386,n5388);
not gate_4889(n5390,n5389);
and gate_4890(n5391,n5086,n5390);
not gate_4891(n5392,n5391);
and gate_4892(n5393,n5384,n5392);
not gate_4893(n5394,n5393);
and gate_4894(po195,n501,n5394);
and gate_4895(n5396,n5277,n5343);
not gate_4896(n5397,n5396);
and gate_4897(n5398,pi255,n5397);
not gate_4898(n5399,n5398);
and gate_4899(n5400,pi208,n5119);
not gate_4900(n5401,n5400);
and gate_4901(n5402,pi209,n5118);
not gate_4902(n5403,n5402);
and gate_4903(n5404,n5401,n5403);
not gate_4904(n5405,n5404);
and gate_4905(n5406,n619,n5405);
not gate_4906(n5407,n5406);
and gate_4907(n5408,n5399,n5407);
not gate_4908(n5409,n5408);
and gate_4909(n5410,n5145,n5409);
not gate_4910(n5411,n5410);
and gate_4911(n5412,pi207,n5144);
not gate_4912(n5413,n5412);
and gate_4913(n5414,n5411,n5413);
not gate_4914(n5415,n5414);
and gate_4915(n5416,n5087,n5415);
not gate_4916(n5417,n5416);
and gate_4917(n5418,pi009,pi048);
not gate_4918(n5419,n5418);
and gate_4919(n5420,n502,pi040);
not gate_4920(n5421,n5420);
and gate_4921(n5422,n5419,n5421);
not gate_4922(n5423,n5422);
and gate_4923(n5424,n5086,n5423);
not gate_4924(n5425,n5424);
and gate_4925(n5426,n5417,n5425);
not gate_4926(n5427,n5426);
and gate_4927(po196,n501,n5427);
and gate_4928(n5429,n5310,n5368);
not gate_4929(n5430,n5429);
and gate_4930(n5431,pi255,n5430);
not gate_4931(n5432,n5431);
and gate_4932(n5433,pi209,n5119);
not gate_4933(n5434,n5433);
and gate_4934(n5435,pi210,n5118);
not gate_4935(n5436,n5435);
and gate_4936(n5437,n5434,n5436);
not gate_4937(n5438,n5437);
and gate_4938(n5439,n619,n5438);
not gate_4939(n5440,n5439);
and gate_4940(n5441,n5432,n5440);
not gate_4941(n5442,n5441);
and gate_4942(n5443,n5145,n5442);
not gate_4943(n5444,n5443);
and gate_4944(n5445,pi208,n5144);
not gate_4945(n5446,n5445);
and gate_4946(n5447,n5444,n5446);
not gate_4947(n5448,n5447);
and gate_4948(n5449,n5087,n5448);
not gate_4949(n5450,n5449);
and gate_4950(n5451,pi009,pi040);
not gate_4951(n5452,n5451);
and gate_4952(n5453,n502,pi032);
not gate_4953(n5454,n5453);
and gate_4954(n5455,n5452,n5454);
not gate_4955(n5456,n5455);
and gate_4956(n5457,n5086,n5456);
not gate_4957(n5458,n5457);
and gate_4958(n5459,n5450,n5458);
not gate_4959(n5460,n5459);
and gate_4960(po197,n501,n5460);
and gate_4961(n5462,n5345,n5401);
not gate_4962(n5463,n5462);
and gate_4963(n5464,pi255,n5463);
not gate_4964(n5465,n5464);
and gate_4965(n5466,pi210,n5119);
not gate_4966(n5467,n5466);
and gate_4967(n5468,pi211,n5118);
not gate_4968(n5469,n5468);
and gate_4969(n5470,n5467,n5469);
not gate_4970(n5471,n5470);
and gate_4971(n5472,n619,n5471);
not gate_4972(n5473,n5472);
and gate_4973(n5474,n5465,n5473);
not gate_4974(n5475,n5474);
and gate_4975(n5476,n5145,n5475);
not gate_4976(n5477,n5476);
and gate_4977(n5478,pi209,n5144);
not gate_4978(n5479,n5478);
and gate_4979(n5480,n5477,n5479);
not gate_4980(n5481,n5480);
and gate_4981(n5482,n5087,n5481);
not gate_4982(n5483,n5482);
and gate_4983(n5484,pi009,pi032);
not gate_4984(n5485,n5484);
and gate_4985(n5486,n502,pi024);
not gate_4986(n5487,n5486);
and gate_4987(n5488,n5485,n5487);
not gate_4988(n5489,n5488);
and gate_4989(n5490,n5086,n5489);
not gate_4990(n5491,n5490);
and gate_4991(n5492,n5483,n5491);
not gate_4992(n5493,n5492);
and gate_4993(po198,n501,n5493);
and gate_4994(n5495,n5370,n5434);
not gate_4995(n5496,n5495);
and gate_4996(n5497,pi255,n5496);
not gate_4997(n5498,n5497);
and gate_4998(n5499,pi211,n5119);
not gate_4999(n5500,n5499);
and gate_5000(n5501,pi212,n5118);
not gate_5001(n5502,n5501);
and gate_5002(n5503,n5500,n5502);
not gate_5003(n5504,n5503);
and gate_5004(n5505,n619,n5504);
not gate_5005(n5506,n5505);
and gate_5006(n5507,n5498,n5506);
not gate_5007(n5508,n5507);
and gate_5008(n5509,n5145,n5508);
not gate_5009(n5510,n5509);
and gate_5010(n5511,pi210,n5144);
not gate_5011(n5512,n5511);
and gate_5012(n5513,n5510,n5512);
not gate_5013(n5514,n5513);
and gate_5014(n5515,n5087,n5514);
not gate_5015(n5516,n5515);
and gate_5016(n5517,pi009,pi024);
not gate_5017(n5518,n5517);
and gate_5018(n5519,n502,pi016);
not gate_5019(n5520,n5519);
and gate_5020(n5521,n5518,n5520);
not gate_5021(n5522,n5521);
and gate_5022(n5523,n5086,n5522);
not gate_5023(n5524,n5523);
and gate_5024(n5525,n5516,n5524);
not gate_5025(n5526,n5525);
and gate_5026(po199,n501,n5526);
and gate_5027(n5528,pi006,n502);
not gate_5028(n5529,n5528);
and gate_5029(n5530,pi009,pi016);
not gate_5030(n5531,n5530);
and gate_5031(n5532,n5529,n5531);
not gate_5032(n5533,n5532);
and gate_5033(n5534,n5086,n5533);
not gate_5034(n5535,n5534);
and gate_5035(n5536,n5403,n5467);
not gate_5036(n5537,n5536);
and gate_5037(n5538,pi255,n5537);
not gate_5038(n5539,n5538);
and gate_5039(n5540,pi213,n5118);
not gate_5040(n5541,n5540);
and gate_5041(n5542,pi212,n5119);
not gate_5042(n5543,n5542);
and gate_5043(n5544,n5541,n5543);
not gate_5044(n5545,n5544);
and gate_5045(n5546,n619,n5545);
not gate_5046(n5547,n5546);
and gate_5047(n5548,n5539,n5547);
not gate_5048(n5549,n5548);
and gate_5049(n5550,n5145,n5549);
not gate_5050(n5551,n5550);
and gate_5051(n5552,pi211,n5144);
not gate_5052(n5553,n5552);
and gate_5053(n5554,n5551,n5553);
not gate_5054(n5555,n5554);
and gate_5055(n5556,n5087,n5555);
not gate_5056(n5557,n5556);
and gate_5057(n5558,n5535,n5557);
not gate_5058(n5559,n5558);
and gate_5059(po200,n501,n5559);
and gate_5060(n5561,pi006,pi009);
not gate_5061(n5562,n5561);
and gate_5062(n5563,n502,pi065);
not gate_5063(n5564,n5563);
and gate_5064(n5565,n5562,n5564);
not gate_5065(n5566,n5565);
and gate_5066(n5567,n5086,n5566);
not gate_5067(n5568,n5567);
and gate_5068(n5569,n5436,n5500);
not gate_5069(n5570,n5569);
and gate_5070(n5571,pi255,n5570);
not gate_5071(n5572,n5571);
and gate_5072(n5573,pi214,n5118);
not gate_5073(n5574,n5573);
and gate_5074(n5575,pi213,n5119);
not gate_5075(n5576,n5575);
and gate_5076(n5577,n5574,n5576);
not gate_5077(n5578,n5577);
and gate_5078(n5579,n619,n5578);
not gate_5079(n5580,n5579);
and gate_5080(n5581,n5572,n5580);
not gate_5081(n5582,n5581);
and gate_5082(n5583,n5145,n5582);
not gate_5083(n5584,n5583);
and gate_5084(n5585,pi212,n5144);
not gate_5085(n5586,n5585);
and gate_5086(n5587,n5584,n5586);
not gate_5087(n5588,n5587);
and gate_5088(n5589,n5087,n5588);
not gate_5089(n5590,n5589);
and gate_5090(n5591,n5568,n5590);
not gate_5091(n5592,n5591);
and gate_5092(po201,n501,n5592);
and gate_5093(n5594,n5469,n5543);
not gate_5094(n5595,n5594);
and gate_5095(n5596,pi255,n5595);
not gate_5096(n5597,n5596);
and gate_5097(n5598,pi214,n5119);
not gate_5098(n5599,n5598);
and gate_5099(n5600,pi215,n5118);
not gate_5100(n5601,n5600);
and gate_5101(n5602,n5599,n5601);
not gate_5102(n5603,n5602);
and gate_5103(n5604,n619,n5603);
not gate_5104(n5605,n5604);
and gate_5105(n5606,n5597,n5605);
not gate_5106(n5607,n5606);
and gate_5107(n5608,n5145,n5607);
not gate_5108(n5609,n5608);
and gate_5109(n5610,pi213,n5144);
not gate_5110(n5611,n5610);
and gate_5111(n5612,n5609,n5611);
not gate_5112(n5613,n5612);
and gate_5113(n5614,n5087,n5613);
not gate_5114(n5615,n5614);
and gate_5115(n5616,pi009,pi065);
not gate_5116(n5617,n5616);
and gate_5117(n5618,n502,pi057);
not gate_5118(n5619,n5618);
and gate_5119(n5620,n5617,n5619);
not gate_5120(n5621,n5620);
and gate_5121(n5622,n5086,n5621);
not gate_5122(n5623,n5622);
and gate_5123(n5624,n5615,n5623);
not gate_5124(n5625,n5624);
and gate_5125(po202,n501,n5625);
and gate_5126(n5627,n502,pi049);
not gate_5127(n5628,n5627);
and gate_5128(n5629,pi009,pi057);
not gate_5129(n5630,n5629);
and gate_5130(n5631,n5628,n5630);
not gate_5131(n5632,n5631);
and gate_5132(n5633,n5086,n5632);
not gate_5133(n5634,n5633);
and gate_5134(n5635,n5502,n5576);
not gate_5135(n5636,n5635);
and gate_5136(n5637,pi255,n5636);
not gate_5137(n5638,n5637);
and gate_5138(n5639,pi215,n5119);
not gate_5139(n5640,n5639);
and gate_5140(n5641,pi216,n5118);
not gate_5141(n5642,n5641);
and gate_5142(n5643,n5640,n5642);
not gate_5143(n5644,n5643);
and gate_5144(n5645,n619,n5644);
not gate_5145(n5646,n5645);
and gate_5146(n5647,n5638,n5646);
not gate_5147(n5648,n5647);
and gate_5148(n5649,n5145,n5648);
not gate_5149(n5650,n5649);
and gate_5150(n5651,pi214,n5144);
not gate_5151(n5652,n5651);
and gate_5152(n5653,n5650,n5652);
not gate_5153(n5654,n5653);
and gate_5154(n5655,n5087,n5654);
not gate_5155(n5656,n5655);
and gate_5156(n5657,n5634,n5656);
not gate_5157(n5658,n5657);
and gate_5158(po203,n501,n5658);
and gate_5159(n5660,pi009,pi049);
not gate_5160(n5661,n5660);
and gate_5161(n5662,n502,pi041);
not gate_5162(n5663,n5662);
and gate_5163(n5664,n5661,n5663);
not gate_5164(n5665,n5664);
and gate_5165(n5666,n5086,n5665);
not gate_5166(n5667,n5666);
and gate_5167(n5668,n5541,n5599);
not gate_5168(n5669,n5668);
and gate_5169(n5670,pi255,n5669);
not gate_5170(n5671,n5670);
and gate_5171(n5672,pi217,n5118);
not gate_5172(n5673,n5672);
and gate_5173(n5674,pi216,n5119);
not gate_5174(n5675,n5674);
and gate_5175(n5676,n5673,n5675);
not gate_5176(n5677,n5676);
and gate_5177(n5678,n619,n5677);
not gate_5178(n5679,n5678);
and gate_5179(n5680,n5671,n5679);
not gate_5180(n5681,n5680);
and gate_5181(n5682,n5145,n5681);
not gate_5182(n5683,n5682);
and gate_5183(n5684,pi215,n5144);
not gate_5184(n5685,n5684);
and gate_5185(n5686,n5683,n5685);
not gate_5186(n5687,n5686);
and gate_5187(n5688,n5087,n5687);
not gate_5188(n5689,n5688);
and gate_5189(n5690,n5667,n5689);
not gate_5190(n5691,n5690);
and gate_5191(po204,n501,n5691);
and gate_5192(n5693,pi009,pi041);
not gate_5193(n5694,n5693);
and gate_5194(n5695,n502,pi033);
not gate_5195(n5696,n5695);
and gate_5196(n5697,n5694,n5696);
not gate_5197(n5698,n5697);
and gate_5198(n5699,n5086,n5698);
not gate_5199(n5700,n5699);
and gate_5200(n5701,n5574,n5640);
not gate_5201(n5702,n5701);
and gate_5202(n5703,pi255,n5702);
not gate_5203(n5704,n5703);
and gate_5204(n5705,pi217,n5119);
not gate_5205(n5706,n5705);
and gate_5206(n5707,pi218,n5118);
not gate_5207(n5708,n5707);
and gate_5208(n5709,n5706,n5708);
not gate_5209(n5710,n5709);
and gate_5210(n5711,n619,n5710);
not gate_5211(n5712,n5711);
and gate_5212(n5713,n5704,n5712);
not gate_5213(n5714,n5713);
and gate_5214(n5715,n5145,n5714);
not gate_5215(n5716,n5715);
and gate_5216(n5717,pi216,n5144);
not gate_5217(n5718,n5717);
and gate_5218(n5719,n5716,n5718);
not gate_5219(n5720,n5719);
and gate_5220(n5721,n5087,n5720);
not gate_5221(n5722,n5721);
and gate_5222(n5723,n5700,n5722);
not gate_5223(n5724,n5723);
and gate_5224(po205,n501,n5724);
and gate_5225(n5726,pi009,pi033);
not gate_5226(n5727,n5726);
and gate_5227(n5728,n502,pi025);
not gate_5228(n5729,n5728);
and gate_5229(n5730,n5727,n5729);
not gate_5230(n5731,n5730);
and gate_5231(n5732,n5086,n5731);
not gate_5232(n5733,n5732);
and gate_5233(n5734,n5601,n5675);
not gate_5234(n5735,n5734);
and gate_5235(n5736,pi255,n5735);
not gate_5236(n5737,n5736);
and gate_5237(n5738,pi218,n5119);
not gate_5238(n5739,n5738);
and gate_5239(n5740,pi219,n5118);
not gate_5240(n5741,n5740);
and gate_5241(n5742,n5739,n5741);
not gate_5242(n5743,n5742);
and gate_5243(n5744,n619,n5743);
not gate_5244(n5745,n5744);
and gate_5245(n5746,n5737,n5745);
not gate_5246(n5747,n5746);
and gate_5247(n5748,n5145,n5747);
not gate_5248(n5749,n5748);
and gate_5249(n5750,pi217,n5144);
not gate_5250(n5751,n5750);
and gate_5251(n5752,n5749,n5751);
not gate_5252(n5753,n5752);
and gate_5253(n5754,n5087,n5753);
not gate_5254(n5755,n5754);
and gate_5255(n5756,n5733,n5755);
not gate_5256(n5757,n5756);
and gate_5257(po206,n501,n5757);
and gate_5258(n5759,pi009,pi025);
not gate_5259(n5760,n5759);
and gate_5260(n5761,n502,pi017);
not gate_5261(n5762,n5761);
and gate_5262(n5763,n5760,n5762);
not gate_5263(n5764,n5763);
and gate_5264(n5765,n5086,n5764);
not gate_5265(n5766,n5765);
and gate_5266(n5767,n5642,n5706);
not gate_5267(n5768,n5767);
and gate_5268(n5769,pi255,n5768);
not gate_5269(n5770,n5769);
and gate_5270(n5771,pi219,n5119);
not gate_5271(n5772,n5771);
and gate_5272(n5773,pi220,n5118);
not gate_5273(n5774,n5773);
and gate_5274(n5775,n5772,n5774);
not gate_5275(n5776,n5775);
and gate_5276(n5777,n619,n5776);
not gate_5277(n5778,n5777);
and gate_5278(n5779,n5770,n5778);
not gate_5279(n5780,n5779);
and gate_5280(n5781,n5145,n5780);
not gate_5281(n5782,n5781);
and gate_5282(n5783,pi218,n5144);
not gate_5283(n5784,n5783);
and gate_5284(n5785,n5782,n5784);
not gate_5285(n5786,n5785);
and gate_5286(n5787,n5087,n5786);
not gate_5287(n5788,n5787);
and gate_5288(n5789,n5766,n5788);
not gate_5289(n5790,n5789);
and gate_5290(po207,n501,n5790);
and gate_5291(n5792,pi007,n502);
not gate_5292(n5793,n5792);
and gate_5293(n5794,pi009,pi017);
not gate_5294(n5795,n5794);
and gate_5295(n5796,n5793,n5795);
not gate_5296(n5797,n5796);
and gate_5297(n5798,n5086,n5797);
not gate_5298(n5799,n5798);
and gate_5299(n5800,n5673,n5739);
not gate_5300(n5801,n5800);
and gate_5301(n5802,pi255,n5801);
not gate_5302(n5803,n5802);
and gate_5303(n5804,pi221,n5118);
not gate_5304(n5805,n5804);
and gate_5305(n5806,pi220,n5119);
not gate_5306(n5807,n5806);
and gate_5307(n5808,n5805,n5807);
not gate_5308(n5809,n5808);
and gate_5309(n5810,n619,n5809);
not gate_5310(n5811,n5810);
and gate_5311(n5812,n5803,n5811);
not gate_5312(n5813,n5812);
and gate_5313(n5814,n5145,n5813);
not gate_5314(n5815,n5814);
and gate_5315(n5816,pi219,n5144);
not gate_5316(n5817,n5816);
and gate_5317(n5818,n5815,n5817);
not gate_5318(n5819,n5818);
and gate_5319(n5820,n5087,n5819);
not gate_5320(n5821,n5820);
and gate_5321(n5822,n5799,n5821);
not gate_5322(n5823,n5822);
and gate_5323(po208,n501,n5823);
and gate_5324(n5825,pi007,pi009);
not gate_5325(n5826,n5825);
and gate_5326(n5827,n502,pi066);
not gate_5327(n5828,n5827);
and gate_5328(n5829,n5826,n5828);
not gate_5329(n5830,n5829);
and gate_5330(n5831,n5086,n5830);
not gate_5331(n5832,n5831);
and gate_5332(n5833,n5708,n5772);
not gate_5333(n5834,n5833);
and gate_5334(n5835,pi255,n5834);
not gate_5335(n5836,n5835);
and gate_5336(n5837,pi222,n5118);
not gate_5337(n5838,n5837);
and gate_5338(n5839,pi221,n5119);
not gate_5339(n5840,n5839);
and gate_5340(n5841,n5838,n5840);
not gate_5341(n5842,n5841);
and gate_5342(n5843,n619,n5842);
not gate_5343(n5844,n5843);
and gate_5344(n5845,n5836,n5844);
not gate_5345(n5846,n5845);
and gate_5346(n5847,n5145,n5846);
not gate_5347(n5848,n5847);
and gate_5348(n5849,pi220,n5144);
not gate_5349(n5850,n5849);
and gate_5350(n5851,n5848,n5850);
not gate_5351(n5852,n5851);
and gate_5352(n5853,n5087,n5852);
not gate_5353(n5854,n5853);
and gate_5354(n5855,n5832,n5854);
not gate_5355(n5856,n5855);
and gate_5356(po209,n501,n5856);
and gate_5357(n5858,n5741,n5807);
not gate_5358(n5859,n5858);
and gate_5359(n5860,pi255,n5859);
not gate_5360(n5861,n5860);
and gate_5361(n5862,pi222,n5119);
not gate_5362(n5863,n5862);
and gate_5363(n5864,pi223,n5118);
not gate_5364(n5865,n5864);
and gate_5365(n5866,n5863,n5865);
not gate_5366(n5867,n5866);
and gate_5367(n5868,n619,n5867);
not gate_5368(n5869,n5868);
and gate_5369(n5870,n5861,n5869);
not gate_5370(n5871,n5870);
and gate_5371(n5872,n5145,n5871);
not gate_5372(n5873,n5872);
and gate_5373(n5874,pi221,n5144);
not gate_5374(n5875,n5874);
and gate_5375(n5876,n5873,n5875);
not gate_5376(n5877,n5876);
and gate_5377(n5878,n5087,n5877);
not gate_5378(n5879,n5878);
and gate_5379(n5880,pi009,pi066);
not gate_5380(n5881,n5880);
and gate_5381(n5882,n502,pi058);
not gate_5382(n5883,n5882);
and gate_5383(n5884,n5881,n5883);
not gate_5384(n5885,n5884);
and gate_5385(n5886,n5086,n5885);
not gate_5386(n5887,n5886);
and gate_5387(n5888,n5879,n5887);
not gate_5388(n5889,n5888);
and gate_5389(po210,n501,n5889);
and gate_5390(n5891,n502,pi050);
not gate_5391(n5892,n5891);
and gate_5392(n5893,pi009,pi058);
not gate_5393(n5894,n5893);
and gate_5394(n5895,n5892,n5894);
not gate_5395(n5896,n5895);
and gate_5396(n5897,n5086,n5896);
not gate_5397(n5898,n5897);
and gate_5398(n5899,n5774,n5840);
not gate_5399(n5900,n5899);
and gate_5400(n5901,pi255,n5900);
not gate_5401(n5902,n5901);
and gate_5402(n5903,pi223,n5119);
not gate_5403(n5904,n5903);
and gate_5404(n5905,pi224,n5118);
not gate_5405(n5906,n5905);
and gate_5406(n5907,n5904,n5906);
not gate_5407(n5908,n5907);
and gate_5408(n5909,n619,n5908);
not gate_5409(n5910,n5909);
and gate_5410(n5911,n5902,n5910);
not gate_5411(n5912,n5911);
and gate_5412(n5913,n5145,n5912);
not gate_5413(n5914,n5913);
and gate_5414(n5915,pi222,n5144);
not gate_5415(n5916,n5915);
and gate_5416(n5917,n5914,n5916);
not gate_5417(n5918,n5917);
and gate_5418(n5919,n5087,n5918);
not gate_5419(n5920,n5919);
and gate_5420(n5921,n5898,n5920);
not gate_5421(n5922,n5921);
and gate_5422(po211,n501,n5922);
and gate_5423(n5924,n5805,n5863);
not gate_5424(n5925,n5924);
and gate_5425(n5926,pi255,n5925);
not gate_5426(n5927,n5926);
and gate_5427(n5928,pi224,n5119);
not gate_5428(n5929,n5928);
and gate_5429(n5930,n5123,n5929);
not gate_5430(n5931,n5930);
and gate_5431(n5932,n619,n5931);
not gate_5432(n5933,n5932);
and gate_5433(n5934,n5927,n5933);
not gate_5434(n5935,n5934);
and gate_5435(n5936,n5145,n5935);
not gate_5436(n5937,n5936);
and gate_5437(n5938,pi223,n5144);
not gate_5438(n5939,n5938);
and gate_5439(n5940,n5937,n5939);
not gate_5440(n5941,n5940);
and gate_5441(n5942,n5087,n5941);
not gate_5442(n5943,n5942);
and gate_5443(n5944,pi009,pi050);
not gate_5444(n5945,n5944);
and gate_5445(n5946,n502,pi042);
not gate_5446(n5947,n5946);
and gate_5447(n5948,n5945,n5947);
not gate_5448(n5949,n5948);
and gate_5449(n5950,n5086,n5949);
not gate_5450(n5951,n5950);
and gate_5451(n5952,n5943,n5951);
not gate_5452(n5953,n5952);
and gate_5453(po212,n501,n5953);
and gate_5454(n5955,n5838,n5904);
not gate_5455(n5956,n5955);
and gate_5456(n5957,pi255,n5956);
not gate_5457(n5958,n5957);
and gate_5458(n5959,pi225,n5119);
not gate_5459(n5960,n5959);
and gate_5460(n5961,n5168,n5960);
not gate_5461(n5962,n5961);
and gate_5462(n5963,n619,n5962);
not gate_5463(n5964,n5963);
and gate_5464(n5965,n5958,n5964);
not gate_5465(n5966,n5965);
and gate_5466(n5967,n5145,n5966);
not gate_5467(n5968,n5967);
and gate_5468(n5969,pi224,n5144);
not gate_5469(n5970,n5969);
and gate_5470(n5971,n5968,n5970);
not gate_5471(n5972,n5971);
and gate_5472(n5973,n5087,n5972);
not gate_5473(n5974,n5973);
and gate_5474(n5975,pi009,pi042);
not gate_5475(n5976,n5975);
and gate_5476(n5977,n502,pi034);
not gate_5477(n5978,n5977);
and gate_5478(n5979,n5976,n5978);
not gate_5479(n5980,n5979);
and gate_5480(n5981,n5086,n5980);
not gate_5481(n5982,n5981);
and gate_5482(n5983,n5974,n5982);
not gate_5483(n5984,n5983);
and gate_5484(po213,n501,n5984);
and gate_5485(n5986,pi009,pi034);
not gate_5486(n5987,n5986);
and gate_5487(n5988,n502,pi026);
not gate_5488(n5989,n5988);
and gate_5489(n5990,n5987,n5989);
not gate_5490(n5991,n5990);
and gate_5491(n5992,n5086,n5991);
not gate_5492(n5993,n5992);
and gate_5493(n5994,pi225,n5144);
not gate_5494(n5995,n5994);
and gate_5495(n5996,n5865,n5929);
not gate_5496(n5997,n5996);
and gate_5497(n5998,pi255,n5997);
not gate_5498(n5999,n5998);
and gate_5499(n6000,n5121,n5195);
not gate_5500(n6001,n6000);
and gate_5501(n6002,n619,n6001);
not gate_5502(n6003,n6002);
and gate_5503(n6004,n5999,n6003);
not gate_5504(n6005,n6004);
and gate_5505(n6006,n5145,n6005);
not gate_5506(n6007,n6006);
and gate_5507(n6008,n5995,n6007);
not gate_5508(n6009,n6008);
and gate_5509(n6010,n5087,n6009);
not gate_5510(n6011,n6010);
and gate_5511(n6012,n5993,n6011);
not gate_5512(n6013,n6012);
and gate_5513(po214,n501,n6013);
and gate_5514(n6015,pi009,pi026);
not gate_5515(n6016,n6015);
and gate_5516(n6017,n502,pi018);
not gate_5517(n6018,n6017);
and gate_5518(n6019,n6016,n6018);
not gate_5519(n6020,n6019);
and gate_5520(n6021,n5086,n6020);
not gate_5521(n6022,n6021);
and gate_5522(n6023,pi226,n5144);
not gate_5523(n6024,n6023);
and gate_5524(n6025,n5166,n5230);
not gate_5525(n6026,n6025);
and gate_5526(n6027,n619,n6026);
not gate_5527(n6028,n6027);
and gate_5528(n6029,n5906,n5960);
not gate_5529(n6030,n6029);
and gate_5530(n6031,pi255,n6030);
not gate_5531(n6032,n6031);
and gate_5532(n6033,n6028,n6032);
not gate_5533(n6034,n6033);
and gate_5534(n6035,n5145,n6034);
not gate_5535(n6036,n6035);
and gate_5536(n6037,n6024,n6036);
not gate_5537(n6038,n6037);
and gate_5538(n6039,n5087,n6038);
not gate_5539(n6040,n6039);
and gate_5540(n6041,n6022,n6040);
not gate_5541(n6042,n6041);
and gate_5542(po215,n501,n6042);
and gate_5543(n6044,pi004,n502);
not gate_5544(n6045,n6044);
and gate_5545(n6046,pi009,pi012);
not gate_5546(n6047,n6046);
and gate_5547(n6048,n6045,n6047);
not gate_5548(n6049,n6048);
and gate_5549(n6050,n5086,n6049);
not gate_5550(n6051,n6050);
and gate_5551(n6052,pi254,n5119);
not gate_5552(n6053,n6052);
and gate_5553(n6054,pi253,n5118);
not gate_5554(n6055,n6054);
and gate_5555(n6056,n6053,n6055);
not gate_5556(n6057,n6056);
and gate_5557(n6058,pi255,n6057);
not gate_5558(n6059,n6058);
and gate_5559(n6060,pi228,n5119);
not gate_5560(n6061,n6060);
and gate_5561(n6062,pi229,n5118);
not gate_5562(n6063,n6062);
and gate_5563(n6064,n6061,n6063);
not gate_5564(n6065,n6064);
and gate_5565(n6066,n619,n6065);
not gate_5566(n6067,n6066);
and gate_5567(n6068,n6059,n6067);
not gate_5568(n6069,n6068);
and gate_5569(n6070,n5145,n6069);
not gate_5570(n6071,n6070);
and gate_5571(n6072,pi227,n5144);
not gate_5572(n6073,n6072);
and gate_5573(n6074,n6071,n6073);
not gate_5574(n6075,n6074);
and gate_5575(n6076,n5087,n6075);
not gate_5576(n6077,n6076);
and gate_5577(n6078,n6051,n6077);
not gate_5578(n6079,n6078);
and gate_5579(po216,n501,n6079);
and gate_5580(n6081,pi004,pi009);
not gate_5581(n6082,n6081);
and gate_5582(n6083,n502,pi063);
not gate_5583(n6084,n6083);
and gate_5584(n6085,n6082,n6084);
not gate_5585(n6086,n6085);
and gate_5586(n6087,n5086,n6086);
not gate_5587(n6088,n6087);
and gate_5588(n6089,pi227,n5119);
not gate_5589(n6090,n6089);
and gate_5590(n6091,pi254,n5118);
not gate_5591(n6092,n6091);
and gate_5592(n6093,n6090,n6092);
not gate_5593(n6094,n6093);
and gate_5594(n6095,pi255,n6094);
not gate_5595(n6096,n6095);
and gate_5596(n6097,pi230,n5118);
not gate_5597(n6098,n6097);
and gate_5598(n6099,pi229,n5119);
not gate_5599(n6100,n6099);
and gate_5600(n6101,n6098,n6100);
not gate_5601(n6102,n6101);
and gate_5602(n6103,n619,n6102);
not gate_5603(n6104,n6103);
and gate_5604(n6105,n6096,n6104);
not gate_5605(n6106,n6105);
and gate_5606(n6107,n5145,n6106);
not gate_5607(n6108,n6107);
and gate_5608(n6109,pi228,n5144);
not gate_5609(n6110,n6109);
and gate_5610(n6111,n6108,n6110);
not gate_5611(n6112,n6111);
and gate_5612(n6113,n5087,n6112);
not gate_5613(n6114,n6113);
and gate_5614(n6115,n6088,n6114);
not gate_5615(n6116,n6115);
and gate_5616(po217,n501,n6116);
and gate_5617(n6118,n502,pi055);
not gate_5618(n6119,n6118);
and gate_5619(n6120,pi009,pi063);
not gate_5620(n6121,n6120);
and gate_5621(n6122,n6119,n6121);
not gate_5622(n6123,n6122);
and gate_5623(n6124,n5086,n6123);
not gate_5624(n6125,n6124);
and gate_5625(n6126,pi227,n5118);
not gate_5626(n6127,n6126);
and gate_5627(n6128,n6061,n6127);
not gate_5628(n6129,n6128);
and gate_5629(n6130,pi255,n6129);
not gate_5630(n6131,n6130);
and gate_5631(n6132,pi230,n5119);
not gate_5632(n6133,n6132);
and gate_5633(n6134,pi231,n5118);
not gate_5634(n6135,n6134);
and gate_5635(n6136,n6133,n6135);
not gate_5636(n6137,n6136);
and gate_5637(n6138,n619,n6137);
not gate_5638(n6139,n6138);
and gate_5639(n6140,n6131,n6139);
not gate_5640(n6141,n6140);
and gate_5641(n6142,n5145,n6141);
not gate_5642(n6143,n6142);
and gate_5643(n6144,pi229,n5144);
not gate_5644(n6145,n6144);
and gate_5645(n6146,n6143,n6145);
not gate_5646(n6147,n6146);
and gate_5647(n6148,n5087,n6147);
not gate_5648(n6149,n6148);
and gate_5649(n6150,n6125,n6149);
not gate_5650(n6151,n6150);
and gate_5651(po218,n501,n6151);
and gate_5652(n6153,pi228,n5118);
not gate_5653(n6154,n6153);
and gate_5654(n6155,n6100,n6154);
not gate_5655(n6156,n6155);
and gate_5656(n6157,pi255,n6156);
not gate_5657(n6158,n6157);
and gate_5658(n6159,pi231,n5119);
not gate_5659(n6160,n6159);
and gate_5660(n6161,pi232,n5118);
not gate_5661(n6162,n6161);
and gate_5662(n6163,n6160,n6162);
not gate_5663(n6164,n6163);
and gate_5664(n6165,n619,n6164);
not gate_5665(n6166,n6165);
and gate_5666(n6167,n6158,n6166);
not gate_5667(n6168,n6167);
and gate_5668(n6169,n5145,n6168);
not gate_5669(n6170,n6169);
and gate_5670(n6171,pi230,n5144);
not gate_5671(n6172,n6171);
and gate_5672(n6173,n6170,n6172);
not gate_5673(n6174,n6173);
and gate_5674(n6175,n5087,n6174);
not gate_5675(n6176,n6175);
and gate_5676(n6177,pi009,pi055);
not gate_5677(n6178,n6177);
and gate_5678(n6179,n502,pi047);
not gate_5679(n6180,n6179);
and gate_5680(n6181,n6178,n6180);
not gate_5681(n6182,n6181);
and gate_5682(n6183,n5086,n6182);
not gate_5683(n6184,n6183);
and gate_5684(n6185,n6176,n6184);
not gate_5685(n6186,n6185);
and gate_5686(po219,n501,n6186);
and gate_5687(n6188,pi003,n502);
not gate_5688(n6189,n6188);
and gate_5689(n6190,pi009,pi047);
not gate_5690(n6191,n6190);
and gate_5691(n6192,n6189,n6191);
not gate_5692(n6193,n6192);
and gate_5693(n6194,n5086,n6193);
not gate_5694(n6195,n6194);
and gate_5695(n6196,n6063,n6133);
not gate_5696(n6197,n6196);
and gate_5697(n6198,pi255,n6197);
not gate_5698(n6199,n6198);
and gate_5699(n6200,pi233,n5118);
not gate_5700(n6201,n6200);
and gate_5701(n6202,pi232,n5119);
not gate_5702(n6203,n6202);
and gate_5703(n6204,n6201,n6203);
not gate_5704(n6205,n6204);
and gate_5705(n6206,n619,n6205);
not gate_5706(n6207,n6206);
and gate_5707(n6208,n6199,n6207);
not gate_5708(n6209,n6208);
and gate_5709(n6210,n5145,n6209);
not gate_5710(n6211,n6210);
and gate_5711(n6212,pi231,n5144);
not gate_5712(n6213,n6212);
and gate_5713(n6214,n6211,n6213);
not gate_5714(n6215,n6214);
and gate_5715(n6216,n5087,n6215);
not gate_5716(n6217,n6216);
and gate_5717(n6218,n6195,n6217);
not gate_5718(n6219,n6218);
and gate_5719(po220,n501,n6219);
and gate_5720(n6221,pi003,pi009);
not gate_5721(n6222,n6221);
and gate_5722(n6223,n502,pi062);
not gate_5723(n6224,n6223);
and gate_5724(n6225,n6222,n6224);
not gate_5725(n6226,n6225);
and gate_5726(n6227,n5086,n6226);
not gate_5727(n6228,n6227);
and gate_5728(n6229,n6098,n6160);
not gate_5729(n6230,n6229);
and gate_5730(n6231,pi255,n6230);
not gate_5731(n6232,n6231);
and gate_5732(n6233,pi234,n5118);
not gate_5733(n6234,n6233);
and gate_5734(n6235,pi233,n5119);
not gate_5735(n6236,n6235);
and gate_5736(n6237,n6234,n6236);
not gate_5737(n6238,n6237);
and gate_5738(n6239,n619,n6238);
not gate_5739(n6240,n6239);
and gate_5740(n6241,n6232,n6240);
not gate_5741(n6242,n6241);
and gate_5742(n6243,n5145,n6242);
not gate_5743(n6244,n6243);
and gate_5744(n6245,pi232,n5144);
not gate_5745(n6246,n6245);
and gate_5746(n6247,n6244,n6246);
not gate_5747(n6248,n6247);
and gate_5748(n6249,n5087,n6248);
not gate_5749(n6250,n6249);
and gate_5750(n6251,n6228,n6250);
not gate_5751(n6252,n6251);
and gate_5752(po221,n501,n6252);
and gate_5753(n6254,n502,pi054);
not gate_5754(n6255,n6254);
and gate_5755(n6256,pi009,pi062);
not gate_5756(n6257,n6256);
and gate_5757(n6258,n6255,n6257);
not gate_5758(n6259,n6258);
and gate_5759(n6260,n5086,n6259);
not gate_5760(n6261,n6260);
and gate_5761(n6262,n6135,n6203);
not gate_5762(n6263,n6262);
and gate_5763(n6264,pi255,n6263);
not gate_5764(n6265,n6264);
and gate_5765(n6266,pi234,n5119);
not gate_5766(n6267,n6266);
and gate_5767(n6268,pi235,n5118);
not gate_5768(n6269,n6268);
and gate_5769(n6270,n6267,n6269);
not gate_5770(n6271,n6270);
and gate_5771(n6272,n619,n6271);
not gate_5772(n6273,n6272);
and gate_5773(n6274,n6265,n6273);
not gate_5774(n6275,n6274);
and gate_5775(n6276,n5145,n6275);
not gate_5776(n6277,n6276);
and gate_5777(n6278,pi233,n5144);
not gate_5778(n6279,n6278);
and gate_5779(n6280,n6277,n6279);
not gate_5780(n6281,n6280);
and gate_5781(n6282,n5087,n6281);
not gate_5782(n6283,n6282);
and gate_5783(n6284,n6261,n6283);
not gate_5784(n6285,n6284);
and gate_5785(po222,n501,n6285);
and gate_5786(n6287,n6162,n6236);
not gate_5787(n6288,n6287);
and gate_5788(n6289,pi255,n6288);
not gate_5789(n6290,n6289);
and gate_5790(n6291,pi235,n5119);
not gate_5791(n6292,n6291);
and gate_5792(n6293,pi236,n5118);
not gate_5793(n6294,n6293);
and gate_5794(n6295,n6292,n6294);
not gate_5795(n6296,n6295);
and gate_5796(n6297,n619,n6296);
not gate_5797(n6298,n6297);
and gate_5798(n6299,n6290,n6298);
not gate_5799(n6300,n6299);
and gate_5800(n6301,n5145,n6300);
not gate_5801(n6302,n6301);
and gate_5802(n6303,pi234,n5144);
not gate_5803(n6304,n6303);
and gate_5804(n6305,n6302,n6304);
not gate_5805(n6306,n6305);
and gate_5806(n6307,n5087,n6306);
not gate_5807(n6308,n6307);
and gate_5808(n6309,pi009,pi054);
not gate_5809(n6310,n6309);
and gate_5810(n6311,n502,pi046);
not gate_5811(n6312,n6311);
and gate_5812(n6313,n6310,n6312);
not gate_5813(n6314,n6313);
and gate_5814(n6315,n5086,n6314);
not gate_5815(n6316,n6315);
and gate_5816(n6317,n6308,n6316);
not gate_5817(n6318,n6317);
and gate_5818(po223,n501,n6318);
and gate_5819(n6320,n6201,n6267);
not gate_5820(n6321,n6320);
and gate_5821(n6322,pi255,n6321);
not gate_5822(n6323,n6322);
and gate_5823(n6324,pi236,n5119);
not gate_5824(n6325,n6324);
and gate_5825(n6326,pi237,n5118);
not gate_5826(n6327,n6326);
and gate_5827(n6328,n6325,n6327);
not gate_5828(n6329,n6328);
and gate_5829(n6330,n619,n6329);
not gate_5830(n6331,n6330);
and gate_5831(n6332,n6323,n6331);
not gate_5832(n6333,n6332);
and gate_5833(n6334,n5145,n6333);
not gate_5834(n6335,n6334);
and gate_5835(n6336,pi235,n5144);
not gate_5836(n6337,n6336);
and gate_5837(n6338,n6335,n6337);
not gate_5838(n6339,n6338);
and gate_5839(n6340,n5087,n6339);
not gate_5840(n6341,n6340);
and gate_5841(n6342,pi009,pi046);
not gate_5842(n6343,n6342);
and gate_5843(n6344,n502,pi038);
not gate_5844(n6345,n6344);
and gate_5845(n6346,n6343,n6345);
not gate_5846(n6347,n6346);
and gate_5847(n6348,n5086,n6347);
not gate_5848(n6349,n6348);
and gate_5849(n6350,n6341,n6349);
not gate_5850(n6351,n6350);
and gate_5851(po224,n501,n6351);
and gate_5852(n6353,n6234,n6292);
not gate_5853(n6354,n6353);
and gate_5854(n6355,pi255,n6354);
not gate_5855(n6356,n6355);
and gate_5856(n6357,pi237,n5119);
not gate_5857(n6358,n6357);
and gate_5858(n6359,pi238,n5118);
not gate_5859(n6360,n6359);
and gate_5860(n6361,n6358,n6360);
not gate_5861(n6362,n6361);
and gate_5862(n6363,n619,n6362);
not gate_5863(n6364,n6363);
and gate_5864(n6365,n6356,n6364);
not gate_5865(n6366,n6365);
and gate_5866(n6367,n5145,n6366);
not gate_5867(n6368,n6367);
and gate_5868(n6369,pi236,n5144);
not gate_5869(n6370,n6369);
and gate_5870(n6371,n6368,n6370);
not gate_5871(n6372,n6371);
and gate_5872(n6373,n5087,n6372);
not gate_5873(n6374,n6373);
and gate_5874(n6375,pi009,pi038);
not gate_5875(n6376,n6375);
and gate_5876(n6377,n502,pi030);
not gate_5877(n6378,n6377);
and gate_5878(n6379,n6376,n6378);
not gate_5879(n6380,n6379);
and gate_5880(n6381,n5086,n6380);
not gate_5881(n6382,n6381);
and gate_5882(n6383,n6374,n6382);
not gate_5883(n6384,n6383);
and gate_5884(po225,n501,n6384);
and gate_5885(n6386,n6269,n6325);
not gate_5886(n6387,n6386);
and gate_5887(n6388,pi255,n6387);
not gate_5888(n6389,n6388);
and gate_5889(n6390,pi238,n5119);
not gate_5890(n6391,n6390);
and gate_5891(n6392,pi239,n5118);
not gate_5892(n6393,n6392);
and gate_5893(n6394,n6391,n6393);
not gate_5894(n6395,n6394);
and gate_5895(n6396,n619,n6395);
not gate_5896(n6397,n6396);
and gate_5897(n6398,n6389,n6397);
not gate_5898(n6399,n6398);
and gate_5899(n6400,n5145,n6399);
not gate_5900(n6401,n6400);
and gate_5901(n6402,pi237,n5144);
not gate_5902(n6403,n6402);
and gate_5903(n6404,n6401,n6403);
not gate_5904(n6405,n6404);
and gate_5905(n6406,n5087,n6405);
not gate_5906(n6407,n6406);
and gate_5907(n6408,pi009,pi030);
not gate_5908(n6409,n6408);
and gate_5909(n6410,n502,pi022);
not gate_5910(n6411,n6410);
and gate_5911(n6412,n6409,n6411);
not gate_5912(n6413,n6412);
and gate_5913(n6414,n5086,n6413);
not gate_5914(n6415,n6414);
and gate_5915(n6416,n6407,n6415);
not gate_5916(n6417,n6416);
and gate_5917(po226,n501,n6417);
and gate_5918(n6419,n6294,n6358);
not gate_5919(n6420,n6419);
and gate_5920(n6421,pi255,n6420);
not gate_5921(n6422,n6421);
and gate_5922(n6423,pi239,n5119);
not gate_5923(n6424,n6423);
and gate_5924(n6425,pi240,n5118);
not gate_5925(n6426,n6425);
and gate_5926(n6427,n6424,n6426);
not gate_5927(n6428,n6427);
and gate_5928(n6429,n619,n6428);
not gate_5929(n6430,n6429);
and gate_5930(n6431,n6422,n6430);
not gate_5931(n6432,n6431);
and gate_5932(n6433,n5145,n6432);
not gate_5933(n6434,n6433);
and gate_5934(n6435,pi238,n5144);
not gate_5935(n6436,n6435);
and gate_5936(n6437,n6434,n6436);
not gate_5937(n6438,n6437);
and gate_5938(n6439,n5087,n6438);
not gate_5939(n6440,n6439);
and gate_5940(n6441,pi009,pi022);
not gate_5941(n6442,n6441);
and gate_5942(n6443,n502,pi014);
not gate_5943(n6444,n6443);
and gate_5944(n6445,n6442,n6444);
not gate_5945(n6446,n6445);
and gate_5946(n6447,n5086,n6446);
not gate_5947(n6448,n6447);
and gate_5948(n6449,n6440,n6448);
not gate_5949(n6450,n6449);
and gate_5950(po227,n501,n6450);
and gate_5951(n6452,pi002,n502);
not gate_5952(n6453,n6452);
and gate_5953(n6454,pi009,pi014);
not gate_5954(n6455,n6454);
and gate_5955(n6456,n6453,n6455);
not gate_5956(n6457,n6456);
and gate_5957(n6458,n5086,n6457);
not gate_5958(n6459,n6458);
and gate_5959(n6460,n6327,n6391);
not gate_5960(n6461,n6460);
and gate_5961(n6462,pi255,n6461);
not gate_5962(n6463,n6462);
and gate_5963(n6464,pi241,n5118);
not gate_5964(n6465,n6464);
and gate_5965(n6466,pi240,n5119);
not gate_5966(n6467,n6466);
and gate_5967(n6468,n6465,n6467);
not gate_5968(n6469,n6468);
and gate_5969(n6470,n619,n6469);
not gate_5970(n6471,n6470);
and gate_5971(n6472,n6463,n6471);
not gate_5972(n6473,n6472);
and gate_5973(n6474,n5145,n6473);
not gate_5974(n6475,n6474);
and gate_5975(n6476,pi239,n5144);
not gate_5976(n6477,n6476);
and gate_5977(n6478,n6475,n6477);
not gate_5978(n6479,n6478);
and gate_5979(n6480,n5087,n6479);
not gate_5980(n6481,n6480);
and gate_5981(n6482,n6459,n6481);
not gate_5982(n6483,n6482);
and gate_5983(po228,n501,n6483);
and gate_5984(n6485,pi002,pi009);
not gate_5985(n6486,n6485);
and gate_5986(n6487,n502,pi061);
not gate_5987(n6488,n6487);
and gate_5988(n6489,n6486,n6488);
not gate_5989(n6490,n6489);
and gate_5990(n6491,n5086,n6490);
not gate_5991(n6492,n6491);
and gate_5992(n6493,n6360,n6424);
not gate_5993(n6494,n6493);
and gate_5994(n6495,pi255,n6494);
not gate_5995(n6496,n6495);
and gate_5996(n6497,pi242,n5118);
not gate_5997(n6498,n6497);
and gate_5998(n6499,pi241,n5119);
not gate_5999(n6500,n6499);
and gate_6000(n6501,n6498,n6500);
not gate_6001(n6502,n6501);
and gate_6002(n6503,n619,n6502);
not gate_6003(n6504,n6503);
and gate_6004(n6505,n6496,n6504);
not gate_6005(n6506,n6505);
and gate_6006(n6507,n5145,n6506);
not gate_6007(n6508,n6507);
and gate_6008(n6509,pi240,n5144);
not gate_6009(n6510,n6509);
and gate_6010(n6511,n6508,n6510);
not gate_6011(n6512,n6511);
and gate_6012(n6513,n5087,n6512);
not gate_6013(n6514,n6513);
and gate_6014(n6515,n6492,n6514);
not gate_6015(n6516,n6515);
and gate_6016(po229,n501,n6516);
and gate_6017(n6518,n502,pi053);
not gate_6018(n6519,n6518);
and gate_6019(n6520,pi009,pi061);
not gate_6020(n6521,n6520);
and gate_6021(n6522,n6519,n6521);
not gate_6022(n6523,n6522);
and gate_6023(n6524,n5086,n6523);
not gate_6024(n6525,n6524);
and gate_6025(n6526,n6393,n6467);
not gate_6026(n6527,n6526);
and gate_6027(n6528,pi255,n6527);
not gate_6028(n6529,n6528);
and gate_6029(n6530,pi242,n5119);
not gate_6030(n6531,n6530);
and gate_6031(n6532,pi243,n5118);
not gate_6032(n6533,n6532);
and gate_6033(n6534,n6531,n6533);
not gate_6034(n6535,n6534);
and gate_6035(n6536,n619,n6535);
not gate_6036(n6537,n6536);
and gate_6037(n6538,n6529,n6537);
not gate_6038(n6539,n6538);
and gate_6039(n6540,n5145,n6539);
not gate_6040(n6541,n6540);
and gate_6041(n6542,pi241,n5144);
not gate_6042(n6543,n6542);
and gate_6043(n6544,n6541,n6543);
not gate_6044(n6545,n6544);
and gate_6045(n6546,n5087,n6545);
not gate_6046(n6547,n6546);
and gate_6047(n6548,n6525,n6547);
not gate_6048(n6549,n6548);
and gate_6049(po230,n501,n6549);
and gate_6050(n6551,n6426,n6500);
not gate_6051(n6552,n6551);
and gate_6052(n6553,pi255,n6552);
not gate_6053(n6554,n6553);
and gate_6054(n6555,pi243,n5119);
not gate_6055(n6556,n6555);
and gate_6056(n6557,pi244,n5118);
not gate_6057(n6558,n6557);
and gate_6058(n6559,n6556,n6558);
not gate_6059(n6560,n6559);
and gate_6060(n6561,n619,n6560);
not gate_6061(n6562,n6561);
and gate_6062(n6563,n6554,n6562);
not gate_6063(n6564,n6563);
and gate_6064(n6565,n5145,n6564);
not gate_6065(n6566,n6565);
and gate_6066(n6567,pi242,n5144);
not gate_6067(n6568,n6567);
and gate_6068(n6569,n6566,n6568);
not gate_6069(n6570,n6569);
and gate_6070(n6571,n5087,n6570);
not gate_6071(n6572,n6571);
and gate_6072(n6573,pi009,pi053);
not gate_6073(n6574,n6573);
and gate_6074(n6575,n502,pi045);
not gate_6075(n6576,n6575);
and gate_6076(n6577,n6574,n6576);
not gate_6077(n6578,n6577);
and gate_6078(n6579,n5086,n6578);
not gate_6079(n6580,n6579);
and gate_6080(n6581,n6572,n6580);
not gate_6081(n6582,n6581);
and gate_6082(po231,n501,n6582);
and gate_6083(n6584,pi009,pi045);
not gate_6084(n6585,n6584);
and gate_6085(n6586,n502,pi037);
not gate_6086(n6587,n6586);
and gate_6087(n6588,n6585,n6587);
not gate_6088(n6589,n6588);
and gate_6089(n6590,n5086,n6589);
not gate_6090(n6591,n6590);
and gate_6091(n6592,n6465,n6531);
not gate_6092(n6593,n6592);
and gate_6093(n6594,pi255,n6593);
not gate_6094(n6595,n6594);
and gate_6095(n6596,pi245,n5118);
not gate_6096(n6597,n6596);
and gate_6097(n6598,pi244,n5119);
not gate_6098(n6599,n6598);
and gate_6099(n6600,n6597,n6599);
not gate_6100(n6601,n6600);
and gate_6101(n6602,n619,n6601);
not gate_6102(n6603,n6602);
and gate_6103(n6604,n6595,n6603);
not gate_6104(n6605,n6604);
and gate_6105(n6606,n5145,n6605);
not gate_6106(n6607,n6606);
and gate_6107(n6608,pi243,n5144);
not gate_6108(n6609,n6608);
and gate_6109(n6610,n6607,n6609);
not gate_6110(n6611,n6610);
and gate_6111(n6612,n5087,n6611);
not gate_6112(n6613,n6612);
and gate_6113(n6614,n6591,n6613);
not gate_6114(n6615,n6614);
and gate_6115(po232,n501,n6615);
and gate_6116(n6617,pi009,pi037);
not gate_6117(n6618,n6617);
and gate_6118(n6619,n502,pi029);
not gate_6119(n6620,n6619);
and gate_6120(n6621,n6618,n6620);
not gate_6121(n6622,n6621);
and gate_6122(n6623,n5086,n6622);
not gate_6123(n6624,n6623);
and gate_6124(n6625,n6498,n6556);
not gate_6125(n6626,n6625);
and gate_6126(n6627,pi255,n6626);
not gate_6127(n6628,n6627);
and gate_6128(n6629,pi245,n5119);
not gate_6129(n6630,n6629);
and gate_6130(n6631,pi246,n5118);
not gate_6131(n6632,n6631);
and gate_6132(n6633,n6630,n6632);
not gate_6133(n6634,n6633);
and gate_6134(n6635,n619,n6634);
not gate_6135(n6636,n6635);
and gate_6136(n6637,n6628,n6636);
not gate_6137(n6638,n6637);
and gate_6138(n6639,n5145,n6638);
not gate_6139(n6640,n6639);
and gate_6140(n6641,pi244,n5144);
not gate_6141(n6642,n6641);
and gate_6142(n6643,n6640,n6642);
not gate_6143(n6644,n6643);
and gate_6144(n6645,n5087,n6644);
not gate_6145(n6646,n6645);
and gate_6146(n6647,n6624,n6646);
not gate_6147(n6648,n6647);
and gate_6148(po233,n501,n6648);
and gate_6149(n6650,pi009,pi029);
not gate_6150(n6651,n6650);
and gate_6151(n6652,n502,pi021);
not gate_6152(n6653,n6652);
and gate_6153(n6654,n6651,n6653);
not gate_6154(n6655,n6654);
and gate_6155(n6656,n5086,n6655);
not gate_6156(n6657,n6656);
and gate_6157(n6658,n6533,n6599);
not gate_6158(n6659,n6658);
and gate_6159(n6660,pi255,n6659);
not gate_6160(n6661,n6660);
and gate_6161(n6662,pi246,n5119);
not gate_6162(n6663,n6662);
and gate_6163(n6664,pi247,n5118);
not gate_6164(n6665,n6664);
and gate_6165(n6666,n6663,n6665);
not gate_6166(n6667,n6666);
and gate_6167(n6668,n619,n6667);
not gate_6168(n6669,n6668);
and gate_6169(n6670,n6661,n6669);
not gate_6170(n6671,n6670);
and gate_6171(n6672,n5145,n6671);
not gate_6172(n6673,n6672);
and gate_6173(n6674,pi245,n5144);
not gate_6174(n6675,n6674);
and gate_6175(n6676,n6673,n6675);
not gate_6176(n6677,n6676);
and gate_6177(n6678,n5087,n6677);
not gate_6178(n6679,n6678);
and gate_6179(n6680,n6657,n6679);
not gate_6180(n6681,n6680);
and gate_6181(po234,n501,n6681);
and gate_6182(n6683,pi009,pi021);
not gate_6183(n6684,n6683);
and gate_6184(n6685,n502,pi013);
not gate_6185(n6686,n6685);
and gate_6186(n6687,n6684,n6686);
not gate_6187(n6688,n6687);
and gate_6188(n6689,n5086,n6688);
not gate_6189(n6690,n6689);
and gate_6190(n6691,n6558,n6630);
not gate_6191(n6692,n6691);
and gate_6192(n6693,pi255,n6692);
not gate_6193(n6694,n6693);
and gate_6194(n6695,pi247,n5119);
not gate_6195(n6696,n6695);
and gate_6196(n6697,pi248,n5118);
not gate_6197(n6698,n6697);
and gate_6198(n6699,n6696,n6698);
not gate_6199(n6700,n6699);
and gate_6200(n6701,n619,n6700);
not gate_6201(n6702,n6701);
and gate_6202(n6703,n6694,n6702);
not gate_6203(n6704,n6703);
and gate_6204(n6705,n5145,n6704);
not gate_6205(n6706,n6705);
and gate_6206(n6707,pi246,n5144);
not gate_6207(n6708,n6707);
and gate_6208(n6709,n6706,n6708);
not gate_6209(n6710,n6709);
and gate_6210(n6711,n5087,n6710);
not gate_6211(n6712,n6711);
and gate_6212(n6713,n6690,n6712);
not gate_6213(n6714,n6713);
and gate_6214(po235,n501,n6714);
and gate_6215(n6716,pi001,n502);
not gate_6216(n6717,n6716);
and gate_6217(n6718,pi009,pi013);
not gate_6218(n6719,n6718);
and gate_6219(n6720,n6717,n6719);
not gate_6220(n6721,n6720);
and gate_6221(n6722,n5086,n6721);
not gate_6222(n6723,n6722);
and gate_6223(n6724,n6597,n6663);
not gate_6224(n6725,n6724);
and gate_6225(n6726,pi255,n6725);
not gate_6226(n6727,n6726);
and gate_6227(n6728,pi249,n5118);
not gate_6228(n6729,n6728);
and gate_6229(n6730,pi248,n5119);
not gate_6230(n6731,n6730);
and gate_6231(n6732,n6729,n6731);
not gate_6232(n6733,n6732);
and gate_6233(n6734,n619,n6733);
not gate_6234(n6735,n6734);
and gate_6235(n6736,n6727,n6735);
not gate_6236(n6737,n6736);
and gate_6237(n6738,n5145,n6737);
not gate_6238(n6739,n6738);
and gate_6239(n6740,pi247,n5144);
not gate_6240(n6741,n6740);
and gate_6241(n6742,n6739,n6741);
not gate_6242(n6743,n6742);
and gate_6243(n6744,n5087,n6743);
not gate_6244(n6745,n6744);
and gate_6245(n6746,n6723,n6745);
not gate_6246(n6747,n6746);
and gate_6247(po236,n501,n6747);
and gate_6248(n6749,pi001,pi009);
not gate_6249(n6750,n6749);
and gate_6250(n6751,n502,pi060);
not gate_6251(n6752,n6751);
and gate_6252(n6753,n6750,n6752);
not gate_6253(n6754,n6753);
and gate_6254(n6755,n5086,n6754);
not gate_6255(n6756,n6755);
and gate_6256(n6757,n6632,n6696);
not gate_6257(n6758,n6757);
and gate_6258(n6759,pi255,n6758);
not gate_6259(n6760,n6759);
and gate_6260(n6761,pi250,n5118);
not gate_6261(n6762,n6761);
and gate_6262(n6763,pi249,n5119);
not gate_6263(n6764,n6763);
and gate_6264(n6765,n6762,n6764);
not gate_6265(n6766,n6765);
and gate_6266(n6767,n619,n6766);
not gate_6267(n6768,n6767);
and gate_6268(n6769,n6760,n6768);
not gate_6269(n6770,n6769);
and gate_6270(n6771,n5145,n6770);
not gate_6271(n6772,n6771);
and gate_6272(n6773,pi248,n5144);
not gate_6273(n6774,n6773);
and gate_6274(n6775,n6772,n6774);
not gate_6275(n6776,n6775);
and gate_6276(n6777,n5087,n6776);
not gate_6277(n6778,n6777);
and gate_6278(n6779,n6756,n6778);
not gate_6279(n6780,n6779);
and gate_6280(po237,n501,n6780);
and gate_6281(n6782,n502,pi052);
not gate_6282(n6783,n6782);
and gate_6283(n6784,pi009,pi060);
not gate_6284(n6785,n6784);
and gate_6285(n6786,n6783,n6785);
not gate_6286(n6787,n6786);
and gate_6287(n6788,n5086,n6787);
not gate_6288(n6789,n6788);
and gate_6289(n6790,n6665,n6731);
not gate_6290(n6791,n6790);
and gate_6291(n6792,pi255,n6791);
not gate_6292(n6793,n6792);
and gate_6293(n6794,pi250,n5119);
not gate_6294(n6795,n6794);
and gate_6295(n6796,pi251,n5118);
not gate_6296(n6797,n6796);
and gate_6297(n6798,n6795,n6797);
not gate_6298(n6799,n6798);
and gate_6299(n6800,n619,n6799);
not gate_6300(n6801,n6800);
and gate_6301(n6802,n6793,n6801);
not gate_6302(n6803,n6802);
and gate_6303(n6804,n5145,n6803);
not gate_6304(n6805,n6804);
and gate_6305(n6806,pi249,n5144);
not gate_6306(n6807,n6806);
and gate_6307(n6808,n6805,n6807);
not gate_6308(n6809,n6808);
and gate_6309(n6810,n5087,n6809);
not gate_6310(n6811,n6810);
and gate_6311(n6812,n6789,n6811);
not gate_6312(n6813,n6812);
and gate_6313(po238,n501,n6813);
and gate_6314(n6815,n6698,n6764);
not gate_6315(n6816,n6815);
and gate_6316(n6817,pi255,n6816);
not gate_6317(n6818,n6817);
and gate_6318(n6819,pi251,n5119);
not gate_6319(n6820,n6819);
and gate_6320(n6821,pi252,n5118);
not gate_6321(n6822,n6821);
and gate_6322(n6823,n6820,n6822);
not gate_6323(n6824,n6823);
and gate_6324(n6825,n619,n6824);
not gate_6325(n6826,n6825);
and gate_6326(n6827,n6818,n6826);
not gate_6327(n6828,n6827);
and gate_6328(n6829,n5145,n6828);
not gate_6329(n6830,n6829);
and gate_6330(n6831,pi250,n5144);
not gate_6331(n6832,n6831);
and gate_6332(n6833,n6830,n6832);
not gate_6333(n6834,n6833);
and gate_6334(n6835,n5087,n6834);
not gate_6335(n6836,n6835);
and gate_6336(n6837,pi009,pi052);
not gate_6337(n6838,n6837);
and gate_6338(n6839,n502,pi044);
not gate_6339(n6840,n6839);
and gate_6340(n6841,n6838,n6840);
not gate_6341(n6842,n6841);
and gate_6342(n6843,n5086,n6842);
not gate_6343(n6844,n6843);
and gate_6344(n6845,n6836,n6844);
not gate_6345(n6846,n6845);
and gate_6346(po239,n501,n6846);
and gate_6347(n6848,n6729,n6795);
not gate_6348(n6849,n6848);
and gate_6349(n6850,pi255,n6849);
not gate_6350(n6851,n6850);
and gate_6351(n6852,pi252,n5119);
not gate_6352(n6853,n6852);
and gate_6353(n6854,n6055,n6853);
not gate_6354(n6855,n6854);
and gate_6355(n6856,n619,n6855);
not gate_6356(n6857,n6856);
and gate_6357(n6858,n6851,n6857);
not gate_6358(n6859,n6858);
and gate_6359(n6860,n5145,n6859);
not gate_6360(n6861,n6860);
and gate_6361(n6862,pi251,n5144);
not gate_6362(n6863,n6862);
and gate_6363(n6864,n6861,n6863);
not gate_6364(n6865,n6864);
and gate_6365(n6866,n5087,n6865);
not gate_6366(n6867,n6866);
and gate_6367(n6868,pi009,pi044);
not gate_6368(n6869,n6868);
and gate_6369(n6870,n502,pi036);
not gate_6370(n6871,n6870);
and gate_6371(n6872,n6869,n6871);
not gate_6372(n6873,n6872);
and gate_6373(n6874,n5086,n6873);
not gate_6374(n6875,n6874);
and gate_6375(n6876,n6867,n6875);
not gate_6376(n6877,n6876);
and gate_6377(po240,n501,n6877);
and gate_6378(n6879,n6762,n6820);
not gate_6379(n6880,n6879);
and gate_6380(n6881,pi255,n6880);
not gate_6381(n6882,n6881);
and gate_6382(n6883,pi253,n5119);
not gate_6383(n6884,n6883);
and gate_6384(n6885,n6092,n6884);
not gate_6385(n6886,n6885);
and gate_6386(n6887,n619,n6886);
not gate_6387(n6888,n6887);
and gate_6388(n6889,n6882,n6888);
not gate_6389(n6890,n6889);
and gate_6390(n6891,n5145,n6890);
not gate_6391(n6892,n6891);
and gate_6392(n6893,pi252,n5144);
not gate_6393(n6894,n6893);
and gate_6394(n6895,n6892,n6894);
not gate_6395(n6896,n6895);
and gate_6396(n6897,n5087,n6896);
not gate_6397(n6898,n6897);
and gate_6398(n6899,pi009,pi036);
not gate_6399(n6900,n6899);
and gate_6400(n6901,n502,pi028);
not gate_6401(n6902,n6901);
and gate_6402(n6903,n6900,n6902);
not gate_6403(n6904,n6903);
and gate_6404(n6905,n5086,n6904);
not gate_6405(n6906,n6905);
and gate_6406(n6907,n6898,n6906);
not gate_6407(n6908,n6907);
and gate_6408(po241,n501,n6908);
and gate_6409(n6910,pi009,pi028);
not gate_6410(n6911,n6910);
and gate_6411(n6912,n502,pi020);
not gate_6412(n6913,n6912);
and gate_6413(n6914,n6911,n6913);
not gate_6414(n6915,n6914);
and gate_6415(n6916,n5086,n6915);
not gate_6416(n6917,n6916);
and gate_6417(n6918,pi253,n5144);
not gate_6418(n6919,n6918);
and gate_6419(n6920,n6797,n6853);
not gate_6420(n6921,n6920);
and gate_6421(n6922,pi255,n6921);
not gate_6422(n6923,n6922);
and gate_6423(n6924,n6053,n6127);
not gate_6424(n6925,n6924);
and gate_6425(n6926,n619,n6925);
not gate_6426(n6927,n6926);
and gate_6427(n6928,n6923,n6927);
not gate_6428(n6929,n6928);
and gate_6429(n6930,n5145,n6929);
not gate_6430(n6931,n6930);
and gate_6431(n6932,n6919,n6931);
not gate_6432(n6933,n6932);
and gate_6433(n6934,n5087,n6933);
not gate_6434(n6935,n6934);
and gate_6435(n6936,n6917,n6935);
not gate_6436(n6937,n6936);
and gate_6437(po242,n501,n6937);
and gate_6438(n6939,pi009,pi020);
not gate_6439(n6940,n6939);
and gate_6440(n6941,n502,pi012);
not gate_6441(n6942,n6941);
and gate_6442(n6943,n6940,n6942);
not gate_6443(n6944,n6943);
and gate_6444(n6945,n5086,n6944);
not gate_6445(n6946,n6945);
and gate_6446(n6947,pi254,n5144);
not gate_6447(n6948,n6947);
and gate_6448(n6949,n6090,n6154);
not gate_6449(n6950,n6949);
and gate_6450(n6951,n619,n6950);
not gate_6451(n6952,n6951);
and gate_6452(n6953,n6822,n6884);
not gate_6453(n6954,n6953);
and gate_6454(n6955,pi255,n6954);
not gate_6455(n6956,n6955);
and gate_6456(n6957,n6952,n6956);
not gate_6457(n6958,n6957);
and gate_6458(n6959,n5145,n6958);
not gate_6459(n6960,n6959);
and gate_6460(n6961,n6948,n6960);
not gate_6461(n6962,n6961);
and gate_6462(n6963,n5087,n6962);
not gate_6463(n6964,n6963);
and gate_6464(n6965,n6946,n6964);
not gate_6465(n6966,n6965);
and gate_6466(po243,n501,n6966);
and gate_6467(n6968,pi255,n630);
not gate_6468(n6969,n6968);
and gate_6469(n6970,pi009,n629);
not gate_6470(n6971,n6970);
and gate_6471(n6972,n6969,n6971);
not gate_6472(po244,n6972);
endmodule
