// Verilog File 
module apex2 (pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
po0,po1,po2);

input pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38;

output po0,po1,po2;

wire n42,n43,n44,n45,n46,n47,n48,n49,n50,
n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,
n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,
n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,
n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,
n91,n92,n93,n94,n95,n96,n97,n98,n99,n100,
n101,n102,n103,n104,n105,n106,n107,n108,n109,n110,
n111,n112,n113,n114,n115,n116,n117,n118,n119,n120,
n121,n122,n123,n124,n125,n126,n127,n128,n129,n130,
n131,n132,n133,n134,n135,n136,n137,n138,n139,n140,
n141,n142,n143,n144,n145,n146,n147,n148,n149,n150,
n151,n152,n153,n154,n155,n156,n157,n158,n159,n160,
n161,n162,n163,n164,n165,n166,n167,n168,n169,n170,
n171,n172,n173,n174,n175,n176,n177,n178,n179,n180,
n181,n182,n183,n184,n185,n186,n187,n188,n189,n190,
n191,n192,n193,n194,n195,n196,n197,n198,n199,n200,
n201,n202,n203,n204,n205,n206,n207,n208,n209,n210,
n211,n212,n213,n214,n215,n216,n217,n218,n219,n220,
n221,n222,n223,n224,n225,n226,n227,n228,n229,n230,
n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,
n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,
n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,
n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,
n271,n272,n273,n274,n275,n276,n277,n278,n279,n280,
n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,
n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,
n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,
n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,
n321,n322,n323,n324,n325,n326,n327,n328,n329,n331,
n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,
n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,
n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,
n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,
n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,
n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,
n392,n393,n394,n395,n396,n397,n398,n399,n400,n401,
n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,
n412,n413,n414,n415,n416,n417,n418,n419,n420,n421,
n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,
n432,n433,n434,n435,n436,n437,n438,n439,n440,n441,
n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,
n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,
n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,
n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,
n482,n483,n484,n485,n486,n487,n488,n490,n491,n492,
n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,
n503,n504,n505,n506,n507,n508,n509,n510,n511,n512,
n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,
n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,
n533,n534,n535,n536,n537,n538,n539,n540,n541,n542,
n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,
n553,n554,n555,n556,n557,n558,n559,n560,n561,n562,
n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,
n573,n574,n575,n576,n577,n578,n579,n580,n581,n582,
n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,
n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,
n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,
n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,
n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,
n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,
n643,n644,n645,n646,n647,n648,n649,n650;
not gate_0(n42,pi00);
not gate_1(n43,pi01);
not gate_2(n44,pi02);
not gate_3(n45,pi04);
not gate_4(n46,pi05);
not gate_5(n47,pi06);
not gate_6(n48,pi07);
not gate_7(n49,pi08);
not gate_8(n50,pi09);
not gate_9(n51,pi10);
not gate_10(n52,pi11);
not gate_11(n53,pi12);
not gate_12(n54,pi13);
not gate_13(n55,pi14);
not gate_14(n56,pi16);
not gate_15(n57,pi17);
not gate_16(n58,pi18);
not gate_17(n59,pi19);
not gate_18(n60,pi20);
not gate_19(n61,pi21);
not gate_20(n62,pi22);
not gate_21(n63,pi23);
not gate_22(n64,pi24);
not gate_23(n65,pi25);
not gate_24(n66,pi26);
not gate_25(n67,pi27);
not gate_26(n68,pi28);
not gate_27(n69,pi29);
not gate_28(n70,pi30);
not gate_29(n71,pi31);
not gate_30(n72,pi32);
not gate_31(n73,pi33);
not gate_32(n74,pi34);
not gate_33(n75,pi35);
and gate_34(n76,pi13,pi14);
not gate_35(n77,n76);
and gate_36(n78,pi12,pi17);
not gate_37(n79,n78);
and gate_38(n80,n64,pi34);
not gate_39(n81,n80);
and gate_40(n82,n74,pi35);
not gate_41(n83,n82);
and gate_42(n84,n81,n83);
not gate_43(n85,n84);
and gate_44(n86,pi20,n61);
not gate_45(n87,n86);
and gate_46(n88,n62,n87);
not gate_47(n89,n88);
and gate_48(n90,pi29,n89);
not gate_49(n91,n90);
and gate_50(n92,pi08,pi32);
not gate_51(n93,n92);
and gate_52(n94,n48,n93);
not gate_53(n95,n94);
and gate_54(n96,n69,n70);
and gate_55(n97,pi36,n96);
and gate_56(n98,n94,n97);
not gate_57(n99,n98);
and gate_58(n100,n91,n99);
and gate_59(n101,n61,pi29);
not gate_60(n102,n101);
and gate_61(n103,n50,pi31);
and gate_62(n104,pi07,n103);
not gate_63(n105,n104);
and gate_64(n106,n102,n104);
not gate_65(n107,n106);
and gate_66(n108,n100,n107);
not gate_67(n109,n108);
and gate_68(n110,n85,n109);
not gate_69(n111,n110);
and gate_70(n112,n42,n60);
not gate_71(n113,n112);
and gate_72(n114,n61,n113);
not gate_73(n115,n114);
and gate_74(n116,n62,n115);
not gate_75(n117,n116);
and gate_76(n118,pi29,n117);
not gate_77(n119,n118);
and gate_78(n120,n105,n119);
and gate_79(n121,n71,n75);
not gate_80(n122,n121);
and gate_81(n123,n49,n121);
not gate_82(n124,n123);
and gate_83(n125,n95,n124);
not gate_84(n126,n125);
and gate_85(n127,n97,n126);
not gate_86(n128,n127);
and gate_87(n129,n120,n128);
not gate_88(n130,n129);
and gate_89(n131,n66,n130);
not gate_90(n132,n131);
and gate_91(n133,pi34,pi36);
and gate_92(n134,n96,n133);
and gate_93(n135,n123,n134);
not gate_94(n136,n135);
and gate_95(n137,n132,n136);
not gate_96(n138,n137);
and gate_97(n139,n64,n138);
not gate_98(n140,n139);
and gate_99(n141,n111,n140);
not gate_100(n142,n141);
and gate_101(n143,n79,n142);
not gate_102(n144,n143);
and gate_103(n145,pi07,n122);
not gate_104(n146,n145);
and gate_105(n147,n61,n70);
and gate_106(n148,n57,n147);
not gate_107(n149,n148);
and gate_108(n150,n43,n57);
not gate_109(n151,n150);
and gate_110(n152,pi12,n151);
not gate_111(n153,n152);
and gate_112(n154,n61,n150);
not gate_113(n155,n154);
and gate_114(n156,pi29,n155);
not gate_115(n157,n156);
and gate_116(n158,n153,n157);
and gate_117(n159,n47,n158);
and gate_118(n160,n45,n46);
and gate_119(n161,n159,n160);
not gate_120(n162,n161);
and gate_121(n163,n149,n162);
not gate_122(n164,n163);
and gate_123(n165,n44,n164);
not gate_124(n166,n165);
and gate_125(n167,n47,pi29);
and gate_126(n168,n160,n167);
not gate_127(n169,n168);
and gate_128(n170,pi30,n169);
not gate_129(n171,n170);
and gate_130(n172,n53,n61);
not gate_131(n173,n172);
and gate_132(n174,n171,n172);
not gate_133(n175,n174);
and gate_134(n176,n166,n175);
not gate_135(n177,n176);
and gate_136(n178,n66,n177);
not gate_137(n179,n178);
and gate_138(n180,n69,pi34);
and gate_139(n181,n153,n180);
and gate_140(n182,n47,n181);
and gate_141(n183,n160,n182);
and gate_142(n184,n44,n183);
not gate_143(n185,n184);
and gate_144(n186,n179,n185);
not gate_145(n187,n186);
and gate_146(n188,n146,n187);
and gate_147(n189,n64,n188);
not gate_148(n190,n189);
and gate_149(n191,n69,n82);
and gate_150(n192,n153,n191);
and gate_151(n193,n48,n192);
and gate_152(n194,n47,n193);
and gate_153(n195,n160,n194);
and gate_154(n196,n44,n195);
not gate_155(n197,n196);
and gate_156(n198,n190,n197);
not gate_157(n199,n198);
and gate_158(n200,n93,n199);
and gate_159(n201,pi36,n200);
not gate_160(n202,n201);
and gate_161(n203,n53,n60);
and gate_162(n204,pi02,n203);
and gate_163(n205,n64,n66);
not gate_164(n206,n205);
and gate_165(n207,n101,n205);
and gate_166(n208,n204,n207);
not gate_167(n209,n208);
and gate_168(n210,n202,n209);
and gate_169(n211,n144,n210);
not gate_170(n212,n211);
and gate_171(n213,n77,n212);
not gate_172(n214,n213);
and gate_173(n215,pi25,pi33);
not gate_174(n216,n215);
and gate_175(n217,pi07,pi31);
not gate_176(n218,n217);
and gate_177(n219,pi10,pi13);
and gate_178(n220,n217,n219);
not gate_179(n221,n220);
and gate_180(n222,n216,n221);
not gate_181(n223,n222);
and gate_182(n224,n55,n223);
not gate_183(n225,n224);
and gate_184(n226,pi14,pi33);
not gate_185(n227,n226);
and gate_186(n228,pi03,n58);
not gate_187(n229,n228);
and gate_188(n230,n52,n59);
not gate_189(n231,n230);
and gate_190(n232,n229,n231);
not gate_191(n233,n232);
and gate_192(n234,pi10,n233);
and gate_193(n235,n217,n234);
not gate_194(n236,n235);
and gate_195(n237,n227,n236);
not gate_196(n238,n237);
and gate_197(n239,n54,n238);
not gate_198(n240,n239);
and gate_199(n241,n225,n240);
not gate_200(n242,n241);
and gate_201(n243,n85,n102);
not gate_202(n244,n243);
and gate_203(n245,n206,n244);
not gate_204(n246,n245);
and gate_205(n247,n242,n246);
not gate_206(n248,n247);
and gate_207(n249,n66,pi29);
and gate_208(n250,n61,n249);
not gate_209(n251,n250);
and gate_210(n252,n44,n180);
not gate_211(n253,n252);
and gate_212(n254,n251,n253);
not gate_213(n255,n254);
and gate_214(n256,pi07,pi35);
not gate_215(n257,n256);
and gate_216(n258,n255,n257);
not gate_217(n259,n258);
and gate_218(n260,n66,n75);
and gate_219(n261,n44,n69);
and gate_220(n262,n260,n261);
not gate_221(n263,n262);
and gate_222(n264,n259,n263);
not gate_223(n265,n264);
and gate_224(n266,n64,n265);
not gate_225(n267,n266);
and gate_226(n268,n44,n48);
and gate_227(n269,n191,n268);
not gate_228(n270,n269);
and gate_229(n271,n267,n270);
not gate_230(n272,n271);
and gate_231(n273,n93,n272);
and gate_232(n274,pi36,n273);
and gate_233(n275,n47,n274);
and gate_234(n276,n160,n275);
not gate_235(n277,n276);
and gate_236(n278,pi02,n64);
and gate_237(n279,n250,n278);
not gate_238(n280,n279);
and gate_239(n281,n277,n280);
not gate_240(n282,n281);
and gate_241(n283,pi10,n232);
not gate_242(n284,n283);
and gate_243(n285,n54,n283);
not gate_244(n286,n285);
and gate_245(n287,n282,n286);
and gate_246(n288,n77,n287);
and gate_247(n289,n50,n288);
and gate_248(n290,n57,n289);
not gate_249(n291,n290);
and gate_250(n292,n248,n291);
not gate_251(n293,n292);
and gate_252(n294,n79,n293);
not gate_253(n295,n294);
and gate_254(n296,n214,n295);
not gate_255(n297,n296);
and gate_256(n298,n67,n297);
and gate_257(n299,n56,n298);
not gate_258(n300,n299);
and gate_259(n301,n71,n72);
and gate_260(n302,n70,n301);
not gate_261(n303,n302);
and gate_262(n304,pi36,n257);
and gate_263(n305,n69,n304);
not gate_264(n306,n305);
and gate_265(n307,n55,n65);
not gate_266(n308,n307);
and gate_267(n309,n102,n308);
and gate_268(n310,pi33,n309);
not gate_269(n311,n310);
and gate_270(n312,n91,n311);
and gate_271(n313,n306,n312);
not gate_272(n314,n313);
and gate_273(n315,n302,n314);
and gate_274(n316,n80,n315);
not gate_275(n317,n316);
and gate_276(n318,n300,n317);
not gate_277(n319,n318);
and gate_278(n320,n63,n319);
not gate_279(n321,n320);
and gate_280(n322,n75,n206);
not gate_281(n323,n322);
and gate_282(n324,n314,n323);
and gate_283(n325,n74,n324);
and gate_284(n326,n302,n325);
not gate_285(n327,n326);
and gate_286(n328,n321,n327);
not gate_287(n329,n328);
and gate_288(po0,n68,n329);
and gate_289(n331,pi17,n173);
not gate_290(n332,n331);
and gate_291(n333,n60,n332);
and gate_292(n334,pi02,n333);
not gate_293(n335,n334);
and gate_294(n336,n61,n62);
not gate_295(n337,n336);
and gate_296(n338,n79,n337);
not gate_297(n339,n338);
and gate_298(n340,n335,n339);
not gate_299(n341,n340);
and gate_300(n342,pi29,n341);
not gate_301(n343,n342);
and gate_302(n344,n216,n218);
not gate_303(n345,n344);
and gate_304(n346,n79,n345);
not gate_305(n347,n346);
and gate_306(n348,n343,n347);
not gate_307(n349,n348);
and gate_308(n350,n66,n349);
not gate_309(n351,n350);
and gate_310(n352,n60,pi29);
not gate_311(n353,n352);
and gate_312(n354,n345,n353);
not gate_313(n355,n354);
and gate_314(n356,pi29,n337);
not gate_315(n357,n356);
and gate_316(n358,n355,n357);
not gate_317(n359,n358);
and gate_318(n360,n79,n359);
and gate_319(n361,pi34,n360);
not gate_320(n362,n361);
and gate_321(n363,n351,n362);
not gate_322(n364,n363);
and gate_323(n365,n64,n364);
not gate_324(n366,n365);
and gate_325(n367,n82,n360);
not gate_326(n368,n367);
and gate_327(n369,n366,n368);
not gate_328(n370,n369);
and gate_329(n371,n77,n370);
not gate_330(n372,n371);
and gate_331(n373,n112,n249);
not gate_332(n374,n373);
and gate_333(n375,n253,n374);
not gate_334(n376,n375);
and gate_335(n377,n54,n73);
not gate_336(n378,n377);
and gate_337(n379,pi14,n378);
not gate_338(n380,n379);
and gate_339(n381,n50,n284);
not gate_340(n382,n381);
and gate_341(n383,pi01,n382);
not gate_342(n384,n383);
and gate_343(n385,n57,n384);
not gate_344(n386,n385);
and gate_345(n387,pi12,n386);
not gate_346(n388,n387);
and gate_347(n389,n380,n388);
not gate_348(n390,n389);
and gate_349(n391,n50,pi13);
and gate_350(n392,n55,n57);
and gate_351(n393,n391,n392);
not gate_352(n394,n393);
and gate_353(n395,n390,n394);
not gate_354(n396,n395);
and gate_355(n397,n376,n396);
and gate_356(n398,n47,n397);
and gate_357(n399,n160,n398);
not gate_358(n400,n399);
and gate_359(n401,n79,n380);
and gate_360(n402,n70,n401);
and gate_361(n403,n66,n402);
and gate_362(n404,n112,n403);
not gate_363(n405,n404);
and gate_364(n406,n400,n405);
not gate_365(n407,n406);
and gate_366(n408,n257,n407);
not gate_367(n409,n408);
and gate_368(n410,n69,n396);
and gate_369(n411,n260,n410);
and gate_370(n412,n47,n411);
and gate_371(n413,n160,n412);
and gate_372(n414,n44,n413);
not gate_373(n415,n414);
and gate_374(n416,n409,n415);
not gate_375(n417,n416);
and gate_376(n418,n64,n417);
not gate_377(n419,n418);
and gate_378(n420,n191,n396);
and gate_379(n421,n48,n420);
and gate_380(n422,n47,n421);
and gate_381(n423,n160,n422);
and gate_382(n424,n44,n423);
not gate_383(n425,n424);
and gate_384(n426,n419,n425);
not gate_385(n427,n426);
and gate_386(n428,n93,n427);
not gate_387(n429,n428);
and gate_388(n430,n48,n49);
not gate_389(n431,n430);
and gate_390(n432,pi31,n72);
not gate_391(n433,n432);
and gate_392(n434,n431,n433);
not gate_393(n435,n434);
and gate_394(n436,n401,n435);
and gate_395(n437,n85,n436);
not gate_396(n438,n437);
and gate_397(n439,pi26,n74);
not gate_398(n440,n439);
and gate_399(n441,n75,n440);
and gate_400(n442,n49,n441);
not gate_401(n443,n442);
and gate_402(n444,n66,n432);
not gate_403(n445,n444);
and gate_404(n446,n443,n445);
not gate_405(n447,n446);
and gate_406(n448,n401,n447);
and gate_407(n449,n64,n448);
not gate_408(n450,n449);
and gate_409(n451,n438,n450);
not gate_410(n452,n451);
and gate_411(n453,n96,n452);
not gate_412(n454,n453);
and gate_413(n455,n429,n454);
not gate_414(n456,n455);
and gate_415(n457,pi37,n456);
not gate_416(n458,n457);
and gate_417(n459,n372,n458);
not gate_418(n460,n459);
and gate_419(n461,n67,n460);
and gate_420(n462,n56,n461);
not gate_421(n463,n462);
and gate_422(n464,n227,n257);
and gate_423(n465,pi37,n464);
not gate_424(n466,n465);
and gate_425(n467,n216,n466);
not gate_426(n468,n467);
and gate_427(n469,n69,n468);
not gate_428(n470,n469);
and gate_429(n471,pi20,n215);
not gate_430(n472,n471);
and gate_431(n473,n357,n472);
and gate_432(n474,n470,n473);
not gate_433(n475,n474);
and gate_434(n476,n302,n475);
and gate_435(n477,n80,n476);
not gate_436(n478,n477);
and gate_437(n479,n463,n478);
not gate_438(n480,n479);
and gate_439(n481,n63,n480);
not gate_440(n482,n481);
and gate_441(n483,n323,n475);
and gate_442(n484,n74,n483);
and gate_443(n485,n302,n484);
not gate_444(n486,n485);
and gate_445(n487,n482,n486);
not gate_446(n488,n487);
and gate_447(po1,n68,n488);
and gate_448(n490,n56,n77);
and gate_449(n491,n67,n79);
and gate_450(n492,n63,n491);
and gate_451(n493,n490,n492);
not gate_452(n494,n493);
and gate_453(n495,n60,n61);
not gate_454(n496,n495);
and gate_455(n497,n493,n495);
not gate_456(n498,n497);
and gate_457(n499,pi29,n498);
not gate_458(n500,n499);
and gate_459(n501,n50,n286);
not gate_460(n502,n501);
and gate_461(n503,pi12,n502);
not gate_462(n504,n503);
and gate_463(n505,pi02,n504);
not gate_464(n506,n505);
and gate_465(n507,pi01,pi12);
not gate_466(n508,n507);
and gate_467(n509,n502,n507);
not gate_468(n510,n509);
and gate_469(n511,n47,n510);
and gate_470(n512,n160,n511);
and gate_471(n513,n44,n512);
not gate_472(n514,n513);
and gate_473(n515,pi30,n514);
not gate_474(n516,n515);
and gate_475(n517,n146,n516);
not gate_476(n518,n517);
and gate_477(n519,n506,n517);
not gate_478(n520,n519);
and gate_479(n521,n54,n232);
not gate_480(n522,n521);
and gate_481(n523,pi10,n522);
not gate_482(n524,n523);
and gate_483(n525,n47,n508);
and gate_484(n526,n160,n525);
and gate_485(n527,n44,n526);
not gate_486(n528,n527);
and gate_487(n529,pi30,n528);
not gate_488(n530,n529);
and gate_489(n531,n75,n530);
and gate_490(n532,n524,n531);
and gate_491(n533,pi09,n532);
not gate_492(n534,n533);
and gate_493(n535,pi02,n53);
not gate_494(n536,n535);
and gate_495(n537,n533,n536);
not gate_496(n538,n537);
and gate_497(n539,n520,n538);
not gate_498(n540,n539);
and gate_499(n541,n93,n540);
and gate_500(n542,n216,n541);
and gate_501(n543,pi38,n542);
not gate_502(n544,n543);
and gate_503(n545,n500,n544);
not gate_504(n546,n545);
and gate_505(n547,n62,n546);
not gate_506(n548,n547);
and gate_507(n549,n518,n534);
not gate_508(n550,n549);
and gate_509(n551,n93,n550);
and gate_510(n552,n216,n551);
and gate_511(n553,pi38,n552);
and gate_512(n554,n69,n553);
not gate_513(n555,n554);
and gate_514(n556,n303,n494);
not gate_515(n557,n556);
and gate_516(n558,n227,n557);
not gate_517(n559,n558);
and gate_518(n560,n555,n558);
and gate_519(n561,n548,n560);
not gate_520(n562,n561);
and gate_521(n563,n66,n562);
not gate_522(n564,n563);
and gate_523(n565,n93,n530);
and gate_524(n566,n232,n565);
and gate_525(n567,n216,n566);
and gate_526(n568,pi38,n567);
and gate_527(n569,n75,n568);
and gate_528(n570,pi09,n569);
not gate_529(n571,n570);
and gate_530(n572,n56,n492);
not gate_531(n573,n572);
and gate_532(n574,n226,n572);
not gate_533(n575,n574);
and gate_534(n576,n571,n575);
not gate_535(n577,n576);
and gate_536(n578,n54,n577);
not gate_537(n579,n578);
and gate_538(n580,n490,n491);
not gate_539(n581,n580);
and gate_540(n582,n303,n581);
not gate_541(n583,n582);
and gate_542(n584,n51,n531);
and gate_543(n585,pi09,n584);
not gate_544(n586,n585);
and gate_545(n587,n518,n586);
not gate_546(n588,n587);
and gate_547(n589,n93,n588);
and gate_548(n590,n216,n589);
and gate_549(n591,pi38,n590);
not gate_550(n592,n591);
and gate_551(n593,n63,n70);
and gate_552(n594,pi14,n593);
and gate_553(n595,pi33,n594);
and gate_554(n596,n301,n595);
not gate_555(n597,n596);
and gate_556(n598,n63,n597);
and gate_557(n599,n592,n598);
and gate_558(n600,n583,n599);
and gate_559(n601,n579,n600);
not gate_560(n602,n601);
and gate_561(n603,n69,n602);
not gate_562(n604,n603);
and gate_563(n605,pi29,n496);
and gate_564(n606,n62,n605);
not gate_565(n607,n606);
and gate_566(n608,n63,n227);
and gate_567(n609,n583,n608);
not gate_568(n610,n609);
and gate_569(n611,pi22,n610);
not gate_570(n612,n611);
and gate_571(n613,n607,n612);
and gate_572(n614,n604,n613);
not gate_573(n615,n614);
and gate_574(n616,pi34,n615);
not gate_575(n617,n616);
and gate_576(n618,n564,n617);
not gate_577(n619,n618);
and gate_578(n620,n64,n619);
not gate_579(n621,n620);
and gate_580(n622,pi13,n303);
not gate_581(n623,n622);
and gate_582(n624,n303,n573);
not gate_583(n625,n624);
and gate_584(n626,pi33,n625);
not gate_585(n627,n626);
and gate_586(n628,n623,n627);
not gate_587(n629,n628);
and gate_588(n630,pi14,n629);
not gate_589(n631,n630);
and gate_590(n632,n93,n516);
and gate_591(n633,n216,n632);
and gate_592(n634,pi38,n633);
and gate_593(n635,n48,n634);
not gate_594(n636,n635);
and gate_595(n637,n625,n636);
and gate_596(n638,n631,n637);
not gate_597(n639,n638);
and gate_598(n640,n69,n639);
not gate_599(n641,n640);
and gate_600(n642,pi22,n559);
not gate_601(n643,n642);
and gate_602(n644,n607,n643);
and gate_603(n645,n641,n644);
not gate_604(n646,n645);
and gate_605(n647,n82,n646);
not gate_606(n648,n647);
and gate_607(n649,n621,n648);
not gate_608(n650,n649);
and gate_609(po2,n68,n650);
endmodule
