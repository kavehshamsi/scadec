// Verilog File 
module i7 (pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,pi133,pi134,pi135,pi136,pi137,pi138,
pi139,pi140,pi141,pi142,pi143,pi144,pi145,pi146,pi147,pi148,
pi149,pi150,pi151,pi152,pi153,pi154,pi155,pi156,pi157,pi158,
pi159,pi160,pi161,pi162,pi163,pi164,pi165,pi166,pi167,pi168,
pi169,pi170,pi171,pi172,pi173,pi174,pi175,pi176,pi177,pi178,
pi179,pi180,pi181,pi182,pi183,pi184,pi185,pi186,pi187,pi188,
pi189,pi190,pi191,pi192,pi193,pi194,pi195,pi196,pi197,pi198,
po00,po01,po02,po03,po04,po05,po06,po07,po08,po09,
po10,po11,po12,po13,po14,po15,po16,po17,po18,po19,
po20,po21,po22,po23,po24,po25,po26,po27,po28,po29,
po30,po31,po32,po33,po34,po35,po36,po37,po38,po39,
po40,po41,po42,po43,po44,po45,po46,po47,po48,po49,
po50,po51,po52,po53,po54,po55,po56,po57,po58,po59,
po60,po61,po62,po63,po64,po65,po66);

input pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,pi133,pi134,pi135,pi136,pi137,pi138,
pi139,pi140,pi141,pi142,pi143,pi144,pi145,pi146,pi147,pi148,
pi149,pi150,pi151,pi152,pi153,pi154,pi155,pi156,pi157,pi158,
pi159,pi160,pi161,pi162,pi163,pi164,pi165,pi166,pi167,pi168,
pi169,pi170,pi171,pi172,pi173,pi174,pi175,pi176,pi177,pi178,
pi179,pi180,pi181,pi182,pi183,pi184,pi185,pi186,pi187,pi188,
pi189,pi190,pi191,pi192,pi193,pi194,pi195,pi196,pi197,pi198;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18,
po19,po20,po21,po22,po23,po24,po25,po26,po27,po28,
po29,po30,po31,po32,po33,po34,po35,po36,po37,po38,
po39,po40,po41,po42,po43,po44,po45,po46,po47,po48,
po49,po50,po51,po52,po53,po54,po55,po56,po57,po58,
po59,po60,po61,po62,po63,po64,po65,po66;

wire n266,n267,n268,n269,n270,n271,n272,n273,n274,
n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,
n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,
n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,
n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,
n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,
n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,
n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,
n345,n346,n347,n348,n349,n351,n352,n353,n354,n355,
n356,n357,n358,n359,n360,n361,n362,n363,n364,n366,
n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,
n377,n378,n379,n381,n382,n383,n384,n385,n386,n387,
n388,n389,n390,n391,n392,n393,n394,n396,n397,n398,
n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,
n409,n411,n412,n413,n414,n415,n416,n417,n418,n419,
n420,n421,n422,n423,n424,n426,n427,n428,n429,n430,
n431,n432,n433,n434,n435,n436,n437,n438,n439,n441,
n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,
n452,n453,n454,n456,n457,n458,n459,n460,n461,n462,
n463,n464,n465,n466,n467,n468,n469,n471,n472,n473,
n474,n475,n476,n477,n478,n479,n480,n481,n482,n483,
n484,n486,n487,n488,n489,n490,n491,n492,n493,n494,
n495,n496,n497,n498,n499,n501,n502,n503,n504,n505,
n506,n507,n508,n509,n510,n511,n512,n513,n514,n516,
n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,
n527,n528,n529,n531,n532,n533,n534,n535,n536,n537,
n538,n539,n540,n541,n542,n543,n544,n546,n547,n548,
n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,
n559,n561,n562,n563,n564,n565,n566,n567,n568,n569,
n570,n571,n572,n573,n574,n576,n577,n578,n579,n580,
n581,n582,n583,n584,n585,n586,n587,n588,n589,n591,
n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,
n602,n603,n604,n606,n607,n608,n609,n610,n611,n612,
n613,n614,n615,n616,n617,n618,n619,n621,n622,n623,
n624,n625,n626,n627,n628,n629,n630,n631,n632,n633,
n634,n636,n637,n638,n639,n640,n641,n642,n643,n644,
n645,n646,n647,n648,n649,n651,n652,n653,n654,n655,
n656,n657,n658,n659,n660,n661,n662,n663,n664,n666,
n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,
n677,n678,n679,n681,n682,n683,n684,n685,n686,n687,
n688,n689,n690,n691,n692,n693,n694,n696,n697,n698,
n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,
n709,n711,n712,n713,n714,n715,n716,n717,n718,n719,
n720,n721,n722,n723,n724,n726,n727,n728,n729,n730,
n731,n732,n733,n734,n735,n736,n737,n738,n739,n741,
n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,
n752,n753,n754,n756,n757,n758,n759,n760,n761,n762,
n763,n764,n765,n766,n767,n768,n769,n770,n771,n772,
n773,n774,n775,n776,n777,n779,n780,n781,n782,n783,
n784,n785,n786,n787,n788,n789,n790,n791,n792,n793,
n794,n795,n796,n797,n798,n799,n800,n802,n803,n804,
n805,n806,n807,n808,n809,n810,n811,n812,n813,n814,
n815,n816,n817,n818,n819,n820,n821,n822,n823,n825,
n826,n827,n828,n829,n830,n831,n832,n833,n834,n835,
n836,n837,n838,n839,n840,n841,n842,n843,n844,n845,
n846,n848,n849,n850,n851,n852,n853,n854,n855,n856,
n857,n858,n859,n860,n861,n862,n863,n864,n865,n866,
n867,n868,n869,n871,n872,n873,n874,n875,n876,n877,
n878,n879,n880,n881,n882,n883,n884,n885,n886,n887,
n888,n889,n890,n891,n892,n894,n895,n896,n897,n898,
n899,n900,n901,n902,n903,n904,n905,n906,n907,n908,
n909,n910,n911,n912,n913,n914,n915,n917,n918,n919,
n920,n921,n922,n923,n924,n925,n926,n927,n928,n929,
n930,n931,n932,n933,n934,n935,n936,n937,n938,n940,
n941,n942,n943,n944,n945,n946,n947,n948,n949,n950,
n951,n952,n953,n954,n955,n956,n957,n958,n959,n960,
n961,n963,n964,n965,n966,n967,n968,n969,n970,n971,
n972,n973,n974,n975,n976,n977,n978,n979,n980,n981,
n982,n983,n984,n986,n987,n988,n989,n990,n991,n992,
n993,n994,n995,n996,n997,n998,n999,n1000,n1001,n1002,
n1003,n1004,n1005,n1006,n1007,n1009,n1010,n1011,n1012,n1013,
n1014,n1015,n1016,n1017,n1018,n1019,n1020,n1021,n1022,n1023,
n1024,n1025,n1026,n1027,n1028,n1029,n1030,n1032,n1033,n1034,
n1035,n1036,n1037,n1038,n1039,n1040,n1041,n1042,n1043,n1044,
n1045,n1046,n1047,n1048,n1049,n1050,n1051,n1052,n1053,n1055,
n1056,n1057,n1058,n1059,n1060,n1061,n1062,n1063,n1064,n1065,
n1066,n1067,n1068,n1069,n1070,n1071,n1072,n1073,n1074,n1075,
n1076,n1078,n1079,n1080,n1081,n1082,n1083,n1084,n1085,n1086,
n1087,n1088,n1089,n1090,n1091,n1092,n1093,n1094,n1095,n1096,
n1097,n1098,n1099,n1101,n1102,n1103,n1104,n1105,n1106,n1107,
n1108,n1109,n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,
n1118,n1119,n1120,n1121,n1122,n1124,n1125,n1126,n1127,n1128,
n1129,n1130,n1131,n1132,n1133,n1134,n1135,n1136,n1137,n1138,
n1139,n1140,n1141,n1142,n1143,n1144,n1145,n1147,n1148,n1149,
n1150,n1151,n1152,n1153,n1154,n1155,n1156,n1157,n1158,n1159,
n1160,n1161,n1162,n1163,n1164,n1165,n1166,n1167,n1168,n1170,
n1171,n1172,n1173,n1174,n1175,n1176,n1177,n1178,n1179,n1180,
n1181,n1182,n1183,n1184,n1185,n1186,n1187,n1188,n1189,n1190,
n1191,n1193,n1194,n1195,n1196,n1197,n1198,n1199,n1200,n1201,
n1202,n1203,n1204,n1205,n1206,n1207,n1208,n1209,n1210,n1211,
n1212,n1213,n1214,n1216,n1217,n1218,n1219,n1220,n1221,n1222,
n1223,n1224,n1225,n1226,n1227,n1228,n1229,n1230,n1231,n1232,
n1233,n1234,n1235,n1236,n1237,n1239,n1240,n1241,n1242,n1243,
n1244,n1245,n1246,n1247,n1248,n1249,n1250,n1251,n1252,n1253,
n1254,n1255,n1256,n1257,n1258,n1259,n1260,n1262,n1263,n1264,
n1265,n1266,n1267,n1268,n1269,n1270,n1271,n1272,n1273,n1274,
n1275,n1276,n1277,n1278,n1279,n1280,n1281,n1282,n1283,n1285,
n1286,n1287,n1288,n1289,n1290,n1291,n1292,n1293,n1294,n1295,
n1296,n1297,n1298,n1299,n1300,n1301,n1302,n1303,n1304,n1305,
n1306,n1308,n1309,n1310,n1311,n1312,n1313,n1314,n1315,n1316,
n1317,n1318,n1319,n1320,n1321,n1322,n1323,n1324,n1325,n1326,
n1327,n1328,n1329,n1331,n1332,n1333,n1334,n1335,n1336,n1337,
n1338,n1339,n1340,n1341,n1342,n1343,n1344,n1345,n1346,n1347,
n1348,n1349,n1350,n1351,n1352,n1354,n1355,n1356,n1357,n1358,
n1359,n1360,n1361,n1362,n1363,n1364,n1365,n1366,n1367,n1368,
n1369,n1370,n1371,n1372,n1373,n1374,n1375,n1377,n1378,n1379,
n1380,n1381,n1382,n1383,n1384,n1385,n1386,n1387,n1388,n1389,
n1390,n1391,n1392,n1393,n1394,n1395,n1396,n1397,n1398,n1400,
n1401,n1402,n1403,n1404,n1405,n1406,n1407,n1408,n1409,n1410,
n1411,n1412,n1413,n1414,n1415,n1416,n1417,n1418,n1419,n1420,
n1421,n1423,n1424,n1425,n1426,n1427,n1428,n1429,n1430,n1431,
n1432,n1433,n1434,n1435,n1436,n1437,n1438,n1439,n1440,n1441,
n1442,n1443,n1444,n1446,n1447,n1448,n1449,n1450,n1451,n1452,
n1453,n1454,n1455,n1456,n1457,n1458,n1459,n1460,n1461,n1462,
n1463,n1464,n1465,n1466,n1467,n1469,n1470,n1471,n1472,n1473,
n1474,n1475,n1476,n1477,n1478,n1479,n1480,n1481,n1482,n1483,
n1484,n1485,n1486,n1487,n1488,n1489,n1490,n1492,n1494,n1495,
n1496,n1497,n1498,n1499,n1500,n1501,n1502,n1503,n1504,n1505,
n1507,n1508,n1509,n1510,n1511,n1512,n1513,n1514,n1515,n1517,
n1518,n1519,n1520,n1521,n1522,n1523,n1524,n1525,n1526,n1527,
n1528,n1529,n1530,n1531,n1532,n1533,n1534,n1536,n1537,n1538,
n1539,n1540,n1541,n1542,n1543,n1544,n1545,n1546,n1547,n1548,
n1549,n1551,n1552,n1553,n1554,n1555,n1556,n1557,n1558,n1559,
n1560,n1561,n1562,n1563,n1564,n1566,n1567,n1568,n1569,n1570,
n1571,n1572,n1573,n1574,n1575,n1576,n1577,n1578,n1579;
not gate_0(n266,pi000);
not gate_1(n267,pi002);
not gate_2(n268,pi058);
not gate_3(n269,pi059);
not gate_4(n270,pi060);
not gate_5(n271,pi061);
not gate_6(n272,pi062);
not gate_7(n273,pi063);
not gate_8(n274,pi064);
not gate_9(n275,pi065);
not gate_10(n276,pi066);
not gate_11(n277,pi067);
not gate_12(n278,pi068);
not gate_13(n279,pi069);
not gate_14(n280,pi070);
not gate_15(n281,pi071);
not gate_16(n282,pi072);
not gate_17(n283,pi073);
not gate_18(n284,pi074);
not gate_19(n285,pi075);
not gate_20(n286,pi076);
not gate_21(n287,pi077);
not gate_22(n288,pi078);
not gate_23(n289,pi079);
not gate_24(n290,pi080);
not gate_25(n291,pi081);
not gate_26(n292,pi082);
not gate_27(n293,pi083);
not gate_28(n294,pi084);
not gate_29(n295,pi085);
not gate_30(n296,pi119);
not gate_31(n297,pi120);
not gate_32(n298,pi121);
not gate_33(n299,pi122);
not gate_34(n300,pi123);
not gate_35(n301,pi124);
not gate_36(n302,pi125);
not gate_37(n303,pi126);
not gate_38(n304,pi127);
not gate_39(n305,pi128);
not gate_40(n306,pi129);
not gate_41(n307,pi130);
not gate_42(n308,pi131);
not gate_43(n309,pi132);
not gate_44(n310,pi133);
not gate_45(n311,pi134);
not gate_46(n312,pi135);
not gate_47(n313,pi136);
not gate_48(n314,pi137);
not gate_49(n315,pi138);
not gate_50(n316,pi139);
not gate_51(n317,pi140);
not gate_52(n318,pi141);
not gate_53(n319,pi142);
not gate_54(n320,pi143);
not gate_55(n321,pi144);
not gate_56(n322,pi145);
not gate_57(n323,pi146);
not gate_58(n324,pi147);
not gate_59(n325,pi148);
not gate_60(n326,pi149);
not gate_61(n327,pi150);
not gate_62(n328,pi184);
not gate_63(n329,pi185);
not gate_64(n330,pi186);
not gate_65(n331,pi187);
not gate_66(n332,pi191);
not gate_67(n333,pi192);
not gate_68(n334,pi193);
not gate_69(n335,pi194);
and gate_70(n336,pi002,n268);
not gate_71(n337,n336);
and gate_72(n338,pi000,n337);
and gate_73(n339,n267,pi030);
not gate_74(n340,n339);
and gate_75(n341,n338,n340);
not gate_76(n342,n341);
and gate_77(n343,pi001,pi002);
not gate_78(n344,n343);
and gate_79(n345,n340,n344);
not gate_80(n346,n345);
and gate_81(n347,n266,n346);
not gate_82(n348,n347);
and gate_83(n349,n342,n348);
not gate_84(po00,n349);
and gate_85(n351,pi002,n269);
not gate_86(n352,n351);
and gate_87(n353,pi000,n352);
and gate_88(n354,n267,pi031);
not gate_89(n355,n354);
and gate_90(n356,n353,n355);
not gate_91(n357,n356);
and gate_92(n358,pi002,pi003);
not gate_93(n359,n358);
and gate_94(n360,n355,n359);
not gate_95(n361,n360);
and gate_96(n362,n266,n361);
not gate_97(n363,n362);
and gate_98(n364,n357,n363);
not gate_99(po01,n364);
and gate_100(n366,pi002,n270);
not gate_101(n367,n366);
and gate_102(n368,pi000,n367);
and gate_103(n369,n267,pi032);
not gate_104(n370,n369);
and gate_105(n371,n368,n370);
not gate_106(n372,n371);
and gate_107(n373,pi002,pi004);
not gate_108(n374,n373);
and gate_109(n375,n370,n374);
not gate_110(n376,n375);
and gate_111(n377,n266,n376);
not gate_112(n378,n377);
and gate_113(n379,n372,n378);
not gate_114(po02,n379);
and gate_115(n381,pi002,n271);
not gate_116(n382,n381);
and gate_117(n383,pi000,n382);
and gate_118(n384,n267,pi033);
not gate_119(n385,n384);
and gate_120(n386,n383,n385);
not gate_121(n387,n386);
and gate_122(n388,pi002,pi005);
not gate_123(n389,n388);
and gate_124(n390,n385,n389);
not gate_125(n391,n390);
and gate_126(n392,n266,n391);
not gate_127(n393,n392);
and gate_128(n394,n387,n393);
not gate_129(po03,n394);
and gate_130(n396,pi002,n272);
not gate_131(n397,n396);
and gate_132(n398,pi000,n397);
and gate_133(n399,n267,pi034);
not gate_134(n400,n399);
and gate_135(n401,n398,n400);
not gate_136(n402,n401);
and gate_137(n403,pi002,pi006);
not gate_138(n404,n403);
and gate_139(n405,n400,n404);
not gate_140(n406,n405);
and gate_141(n407,n266,n406);
not gate_142(n408,n407);
and gate_143(n409,n402,n408);
not gate_144(po04,n409);
and gate_145(n411,pi002,n273);
not gate_146(n412,n411);
and gate_147(n413,pi000,n412);
and gate_148(n414,n267,pi035);
not gate_149(n415,n414);
and gate_150(n416,n413,n415);
not gate_151(n417,n416);
and gate_152(n418,pi002,pi007);
not gate_153(n419,n418);
and gate_154(n420,n415,n419);
not gate_155(n421,n420);
and gate_156(n422,n266,n421);
not gate_157(n423,n422);
and gate_158(n424,n417,n423);
not gate_159(po05,n424);
and gate_160(n426,pi002,n274);
not gate_161(n427,n426);
and gate_162(n428,pi000,n427);
and gate_163(n429,n267,pi036);
not gate_164(n430,n429);
and gate_165(n431,n428,n430);
not gate_166(n432,n431);
and gate_167(n433,pi002,pi008);
not gate_168(n434,n433);
and gate_169(n435,n430,n434);
not gate_170(n436,n435);
and gate_171(n437,n266,n436);
not gate_172(n438,n437);
and gate_173(n439,n432,n438);
not gate_174(po06,n439);
and gate_175(n441,pi002,n275);
not gate_176(n442,n441);
and gate_177(n443,pi000,n442);
and gate_178(n444,n267,pi037);
not gate_179(n445,n444);
and gate_180(n446,n443,n445);
not gate_181(n447,n446);
and gate_182(n448,pi002,pi009);
not gate_183(n449,n448);
and gate_184(n450,n445,n449);
not gate_185(n451,n450);
and gate_186(n452,n266,n451);
not gate_187(n453,n452);
and gate_188(n454,n447,n453);
not gate_189(po07,n454);
and gate_190(n456,pi002,n276);
not gate_191(n457,n456);
and gate_192(n458,pi000,n457);
and gate_193(n459,n267,pi038);
not gate_194(n460,n459);
and gate_195(n461,n458,n460);
not gate_196(n462,n461);
and gate_197(n463,pi002,pi010);
not gate_198(n464,n463);
and gate_199(n465,n460,n464);
not gate_200(n466,n465);
and gate_201(n467,n266,n466);
not gate_202(n468,n467);
and gate_203(n469,n462,n468);
not gate_204(po08,n469);
and gate_205(n471,pi002,n277);
not gate_206(n472,n471);
and gate_207(n473,pi000,n472);
and gate_208(n474,n267,pi039);
not gate_209(n475,n474);
and gate_210(n476,n473,n475);
not gate_211(n477,n476);
and gate_212(n478,pi002,pi011);
not gate_213(n479,n478);
and gate_214(n480,n475,n479);
not gate_215(n481,n480);
and gate_216(n482,n266,n481);
not gate_217(n483,n482);
and gate_218(n484,n477,n483);
not gate_219(po09,n484);
and gate_220(n486,pi002,n278);
not gate_221(n487,n486);
and gate_222(n488,pi000,n487);
and gate_223(n489,n267,pi040);
not gate_224(n490,n489);
and gate_225(n491,n488,n490);
not gate_226(n492,n491);
and gate_227(n493,pi002,pi012);
not gate_228(n494,n493);
and gate_229(n495,n490,n494);
not gate_230(n496,n495);
and gate_231(n497,n266,n496);
not gate_232(n498,n497);
and gate_233(n499,n492,n498);
not gate_234(po10,n499);
and gate_235(n501,pi002,n279);
not gate_236(n502,n501);
and gate_237(n503,pi000,n502);
and gate_238(n504,n267,pi041);
not gate_239(n505,n504);
and gate_240(n506,n503,n505);
not gate_241(n507,n506);
and gate_242(n508,pi002,pi013);
not gate_243(n509,n508);
and gate_244(n510,n505,n509);
not gate_245(n511,n510);
and gate_246(n512,n266,n511);
not gate_247(n513,n512);
and gate_248(n514,n507,n513);
not gate_249(po11,n514);
and gate_250(n516,pi002,n280);
not gate_251(n517,n516);
and gate_252(n518,pi000,n517);
and gate_253(n519,n267,pi042);
not gate_254(n520,n519);
and gate_255(n521,n518,n520);
not gate_256(n522,n521);
and gate_257(n523,pi002,pi014);
not gate_258(n524,n523);
and gate_259(n525,n520,n524);
not gate_260(n526,n525);
and gate_261(n527,n266,n526);
not gate_262(n528,n527);
and gate_263(n529,n522,n528);
not gate_264(po12,n529);
and gate_265(n531,pi002,n281);
not gate_266(n532,n531);
and gate_267(n533,pi000,n532);
and gate_268(n534,n267,pi043);
not gate_269(n535,n534);
and gate_270(n536,n533,n535);
not gate_271(n537,n536);
and gate_272(n538,pi002,pi015);
not gate_273(n539,n538);
and gate_274(n540,n535,n539);
not gate_275(n541,n540);
and gate_276(n542,n266,n541);
not gate_277(n543,n542);
and gate_278(n544,n537,n543);
not gate_279(po13,n544);
and gate_280(n546,pi002,n282);
not gate_281(n547,n546);
and gate_282(n548,pi000,n547);
and gate_283(n549,n267,pi044);
not gate_284(n550,n549);
and gate_285(n551,n548,n550);
not gate_286(n552,n551);
and gate_287(n553,pi002,pi016);
not gate_288(n554,n553);
and gate_289(n555,n550,n554);
not gate_290(n556,n555);
and gate_291(n557,n266,n556);
not gate_292(n558,n557);
and gate_293(n559,n552,n558);
not gate_294(po14,n559);
and gate_295(n561,pi002,n283);
not gate_296(n562,n561);
and gate_297(n563,pi000,n562);
and gate_298(n564,n267,pi045);
not gate_299(n565,n564);
and gate_300(n566,n563,n565);
not gate_301(n567,n566);
and gate_302(n568,pi002,pi017);
not gate_303(n569,n568);
and gate_304(n570,n565,n569);
not gate_305(n571,n570);
and gate_306(n572,n266,n571);
not gate_307(n573,n572);
and gate_308(n574,n567,n573);
not gate_309(po15,n574);
and gate_310(n576,pi002,n284);
not gate_311(n577,n576);
and gate_312(n578,pi000,n577);
and gate_313(n579,n267,pi046);
not gate_314(n580,n579);
and gate_315(n581,n578,n580);
not gate_316(n582,n581);
and gate_317(n583,pi002,pi018);
not gate_318(n584,n583);
and gate_319(n585,n580,n584);
not gate_320(n586,n585);
and gate_321(n587,n266,n586);
not gate_322(n588,n587);
and gate_323(n589,n582,n588);
not gate_324(po16,n589);
and gate_325(n591,pi002,n285);
not gate_326(n592,n591);
and gate_327(n593,pi000,n592);
and gate_328(n594,n267,pi047);
not gate_329(n595,n594);
and gate_330(n596,n593,n595);
not gate_331(n597,n596);
and gate_332(n598,pi002,pi019);
not gate_333(n599,n598);
and gate_334(n600,n595,n599);
not gate_335(n601,n600);
and gate_336(n602,n266,n601);
not gate_337(n603,n602);
and gate_338(n604,n597,n603);
not gate_339(po17,n604);
and gate_340(n606,pi002,n286);
not gate_341(n607,n606);
and gate_342(n608,pi000,n607);
and gate_343(n609,n267,pi048);
not gate_344(n610,n609);
and gate_345(n611,n608,n610);
not gate_346(n612,n611);
and gate_347(n613,pi002,pi020);
not gate_348(n614,n613);
and gate_349(n615,n610,n614);
not gate_350(n616,n615);
and gate_351(n617,n266,n616);
not gate_352(n618,n617);
and gate_353(n619,n612,n618);
not gate_354(po18,n619);
and gate_355(n621,pi002,n287);
not gate_356(n622,n621);
and gate_357(n623,pi000,n622);
and gate_358(n624,n267,pi049);
not gate_359(n625,n624);
and gate_360(n626,n623,n625);
not gate_361(n627,n626);
and gate_362(n628,pi002,pi021);
not gate_363(n629,n628);
and gate_364(n630,n625,n629);
not gate_365(n631,n630);
and gate_366(n632,n266,n631);
not gate_367(n633,n632);
and gate_368(n634,n627,n633);
not gate_369(po19,n634);
and gate_370(n636,pi002,n288);
not gate_371(n637,n636);
and gate_372(n638,pi000,n637);
and gate_373(n639,n267,pi050);
not gate_374(n640,n639);
and gate_375(n641,n638,n640);
not gate_376(n642,n641);
and gate_377(n643,pi002,pi022);
not gate_378(n644,n643);
and gate_379(n645,n640,n644);
not gate_380(n646,n645);
and gate_381(n647,n266,n646);
not gate_382(n648,n647);
and gate_383(n649,n642,n648);
not gate_384(po20,n649);
and gate_385(n651,pi002,n289);
not gate_386(n652,n651);
and gate_387(n653,pi000,n652);
and gate_388(n654,n267,pi051);
not gate_389(n655,n654);
and gate_390(n656,n653,n655);
not gate_391(n657,n656);
and gate_392(n658,pi002,pi023);
not gate_393(n659,n658);
and gate_394(n660,n655,n659);
not gate_395(n661,n660);
and gate_396(n662,n266,n661);
not gate_397(n663,n662);
and gate_398(n664,n657,n663);
not gate_399(po21,n664);
and gate_400(n666,pi002,n290);
not gate_401(n667,n666);
and gate_402(n668,pi000,n667);
and gate_403(n669,n267,pi052);
not gate_404(n670,n669);
and gate_405(n671,n668,n670);
not gate_406(n672,n671);
and gate_407(n673,pi002,pi024);
not gate_408(n674,n673);
and gate_409(n675,n670,n674);
not gate_410(n676,n675);
and gate_411(n677,n266,n676);
not gate_412(n678,n677);
and gate_413(n679,n672,n678);
not gate_414(po22,n679);
and gate_415(n681,pi002,n291);
not gate_416(n682,n681);
and gate_417(n683,pi000,n682);
and gate_418(n684,n267,pi053);
not gate_419(n685,n684);
and gate_420(n686,n683,n685);
not gate_421(n687,n686);
and gate_422(n688,pi002,pi025);
not gate_423(n689,n688);
and gate_424(n690,n685,n689);
not gate_425(n691,n690);
and gate_426(n692,n266,n691);
not gate_427(n693,n692);
and gate_428(n694,n687,n693);
not gate_429(po23,n694);
and gate_430(n696,pi002,n292);
not gate_431(n697,n696);
and gate_432(n698,pi000,n697);
and gate_433(n699,n267,pi054);
not gate_434(n700,n699);
and gate_435(n701,n698,n700);
not gate_436(n702,n701);
and gate_437(n703,pi002,pi026);
not gate_438(n704,n703);
and gate_439(n705,n700,n704);
not gate_440(n706,n705);
and gate_441(n707,n266,n706);
not gate_442(n708,n707);
and gate_443(n709,n702,n708);
not gate_444(po24,n709);
and gate_445(n711,pi002,n293);
not gate_446(n712,n711);
and gate_447(n713,pi000,n712);
and gate_448(n714,n267,pi055);
not gate_449(n715,n714);
and gate_450(n716,n713,n715);
not gate_451(n717,n716);
and gate_452(n718,pi002,pi027);
not gate_453(n719,n718);
and gate_454(n720,n715,n719);
not gate_455(n721,n720);
and gate_456(n722,n266,n721);
not gate_457(n723,n722);
and gate_458(n724,n717,n723);
not gate_459(po25,n724);
and gate_460(n726,pi002,n294);
not gate_461(n727,n726);
and gate_462(n728,pi000,n727);
and gate_463(n729,n267,pi056);
not gate_464(n730,n729);
and gate_465(n731,n728,n730);
not gate_466(n732,n731);
and gate_467(n733,pi002,pi028);
not gate_468(n734,n733);
and gate_469(n735,n730,n734);
not gate_470(n736,n735);
and gate_471(n737,n266,n736);
not gate_472(n738,n737);
and gate_473(n739,n732,n738);
not gate_474(po26,n739);
and gate_475(n741,pi002,n295);
not gate_476(n742,n741);
and gate_477(n743,pi000,n742);
and gate_478(n744,n267,pi057);
not gate_479(n745,n744);
and gate_480(n746,n743,n745);
not gate_481(n747,n746);
and gate_482(n748,pi002,pi029);
not gate_483(n749,n748);
and gate_484(n750,n745,n749);
not gate_485(n751,n750);
and gate_486(n752,n266,n751);
not gate_487(n753,n752);
and gate_488(n754,n747,n753);
not gate_489(po27,n754);
and gate_490(n756,n267,n296);
not gate_491(n757,n756);
and gate_492(n758,pi087,n757);
not gate_493(n759,n758);
and gate_494(n760,pi000,n759);
not gate_495(n761,n760);
and gate_496(n762,pi002,pi151);
and gate_497(n763,pi000,n762);
not gate_498(n764,n763);
and gate_499(n765,pi002,pi086);
not gate_500(n766,n765);
and gate_501(n767,n267,pi119);
not gate_502(n768,n767);
and gate_503(n769,n766,n768);
not gate_504(n770,n769);
and gate_505(n771,n266,n770);
not gate_506(n772,n771);
and gate_507(n773,n764,n772);
not gate_508(n774,n773);
and gate_509(n775,pi087,n774);
not gate_510(n776,n775);
and gate_511(n777,n761,n776);
not gate_512(po28,n777);
and gate_513(n779,n267,n297);
not gate_514(n780,n779);
and gate_515(n781,pi087,n780);
not gate_516(n782,n781);
and gate_517(n783,pi000,n782);
not gate_518(n784,n783);
and gate_519(n785,pi002,pi152);
and gate_520(n786,pi000,n785);
not gate_521(n787,n786);
and gate_522(n788,pi002,pi088);
not gate_523(n789,n788);
and gate_524(n790,n267,pi120);
not gate_525(n791,n790);
and gate_526(n792,n789,n791);
not gate_527(n793,n792);
and gate_528(n794,n266,n793);
not gate_529(n795,n794);
and gate_530(n796,n787,n795);
not gate_531(n797,n796);
and gate_532(n798,pi087,n797);
not gate_533(n799,n798);
and gate_534(n800,n784,n799);
not gate_535(po29,n800);
and gate_536(n802,n267,n298);
not gate_537(n803,n802);
and gate_538(n804,pi087,n803);
not gate_539(n805,n804);
and gate_540(n806,pi000,n805);
not gate_541(n807,n806);
and gate_542(n808,pi002,pi153);
and gate_543(n809,pi000,n808);
not gate_544(n810,n809);
and gate_545(n811,pi002,pi089);
not gate_546(n812,n811);
and gate_547(n813,n267,pi121);
not gate_548(n814,n813);
and gate_549(n815,n812,n814);
not gate_550(n816,n815);
and gate_551(n817,n266,n816);
not gate_552(n818,n817);
and gate_553(n819,n810,n818);
not gate_554(n820,n819);
and gate_555(n821,pi087,n820);
not gate_556(n822,n821);
and gate_557(n823,n807,n822);
not gate_558(po30,n823);
and gate_559(n825,n267,n299);
not gate_560(n826,n825);
and gate_561(n827,pi087,n826);
not gate_562(n828,n827);
and gate_563(n829,pi000,n828);
not gate_564(n830,n829);
and gate_565(n831,pi002,pi154);
and gate_566(n832,pi000,n831);
not gate_567(n833,n832);
and gate_568(n834,pi002,pi090);
not gate_569(n835,n834);
and gate_570(n836,n267,pi122);
not gate_571(n837,n836);
and gate_572(n838,n835,n837);
not gate_573(n839,n838);
and gate_574(n840,n266,n839);
not gate_575(n841,n840);
and gate_576(n842,n833,n841);
not gate_577(n843,n842);
and gate_578(n844,pi087,n843);
not gate_579(n845,n844);
and gate_580(n846,n830,n845);
not gate_581(po31,n846);
and gate_582(n848,n267,n300);
not gate_583(n849,n848);
and gate_584(n850,pi087,n849);
not gate_585(n851,n850);
and gate_586(n852,pi000,n851);
not gate_587(n853,n852);
and gate_588(n854,pi002,pi155);
and gate_589(n855,pi000,n854);
not gate_590(n856,n855);
and gate_591(n857,pi002,pi091);
not gate_592(n858,n857);
and gate_593(n859,n267,pi123);
not gate_594(n860,n859);
and gate_595(n861,n858,n860);
not gate_596(n862,n861);
and gate_597(n863,n266,n862);
not gate_598(n864,n863);
and gate_599(n865,n856,n864);
not gate_600(n866,n865);
and gate_601(n867,pi087,n866);
not gate_602(n868,n867);
and gate_603(n869,n853,n868);
not gate_604(po32,n869);
and gate_605(n871,n267,n301);
not gate_606(n872,n871);
and gate_607(n873,pi087,n872);
not gate_608(n874,n873);
and gate_609(n875,pi000,n874);
not gate_610(n876,n875);
and gate_611(n877,pi002,pi156);
and gate_612(n878,pi000,n877);
not gate_613(n879,n878);
and gate_614(n880,pi002,pi092);
not gate_615(n881,n880);
and gate_616(n882,n267,pi124);
not gate_617(n883,n882);
and gate_618(n884,n881,n883);
not gate_619(n885,n884);
and gate_620(n886,n266,n885);
not gate_621(n887,n886);
and gate_622(n888,n879,n887);
not gate_623(n889,n888);
and gate_624(n890,pi087,n889);
not gate_625(n891,n890);
and gate_626(n892,n876,n891);
not gate_627(po33,n892);
and gate_628(n894,n267,n302);
not gate_629(n895,n894);
and gate_630(n896,pi087,n895);
not gate_631(n897,n896);
and gate_632(n898,pi000,n897);
not gate_633(n899,n898);
and gate_634(n900,pi002,pi157);
and gate_635(n901,pi000,n900);
not gate_636(n902,n901);
and gate_637(n903,pi002,pi093);
not gate_638(n904,n903);
and gate_639(n905,n267,pi125);
not gate_640(n906,n905);
and gate_641(n907,n904,n906);
not gate_642(n908,n907);
and gate_643(n909,n266,n908);
not gate_644(n910,n909);
and gate_645(n911,n902,n910);
not gate_646(n912,n911);
and gate_647(n913,pi087,n912);
not gate_648(n914,n913);
and gate_649(n915,n899,n914);
not gate_650(po34,n915);
and gate_651(n917,n267,n303);
not gate_652(n918,n917);
and gate_653(n919,pi087,n918);
not gate_654(n920,n919);
and gate_655(n921,pi000,n920);
not gate_656(n922,n921);
and gate_657(n923,pi002,pi158);
and gate_658(n924,pi000,n923);
not gate_659(n925,n924);
and gate_660(n926,pi002,pi094);
not gate_661(n927,n926);
and gate_662(n928,n267,pi126);
not gate_663(n929,n928);
and gate_664(n930,n927,n929);
not gate_665(n931,n930);
and gate_666(n932,n266,n931);
not gate_667(n933,n932);
and gate_668(n934,n925,n933);
not gate_669(n935,n934);
and gate_670(n936,pi087,n935);
not gate_671(n937,n936);
and gate_672(n938,n922,n937);
not gate_673(po35,n938);
and gate_674(n940,n267,n304);
not gate_675(n941,n940);
and gate_676(n942,pi087,n941);
not gate_677(n943,n942);
and gate_678(n944,pi000,n943);
not gate_679(n945,n944);
and gate_680(n946,pi002,pi159);
and gate_681(n947,pi000,n946);
not gate_682(n948,n947);
and gate_683(n949,pi002,pi095);
not gate_684(n950,n949);
and gate_685(n951,n267,pi127);
not gate_686(n952,n951);
and gate_687(n953,n950,n952);
not gate_688(n954,n953);
and gate_689(n955,n266,n954);
not gate_690(n956,n955);
and gate_691(n957,n948,n956);
not gate_692(n958,n957);
and gate_693(n959,pi087,n958);
not gate_694(n960,n959);
and gate_695(n961,n945,n960);
not gate_696(po36,n961);
and gate_697(n963,n267,n305);
not gate_698(n964,n963);
and gate_699(n965,pi087,n964);
not gate_700(n966,n965);
and gate_701(n967,pi000,n966);
not gate_702(n968,n967);
and gate_703(n969,pi002,pi160);
and gate_704(n970,pi000,n969);
not gate_705(n971,n970);
and gate_706(n972,pi002,pi096);
not gate_707(n973,n972);
and gate_708(n974,n267,pi128);
not gate_709(n975,n974);
and gate_710(n976,n973,n975);
not gate_711(n977,n976);
and gate_712(n978,n266,n977);
not gate_713(n979,n978);
and gate_714(n980,n971,n979);
not gate_715(n981,n980);
and gate_716(n982,pi087,n981);
not gate_717(n983,n982);
and gate_718(n984,n968,n983);
not gate_719(po37,n984);
and gate_720(n986,n267,n306);
not gate_721(n987,n986);
and gate_722(n988,pi087,n987);
not gate_723(n989,n988);
and gate_724(n990,pi000,n989);
not gate_725(n991,n990);
and gate_726(n992,pi002,pi161);
and gate_727(n993,pi000,n992);
not gate_728(n994,n993);
and gate_729(n995,pi002,pi097);
not gate_730(n996,n995);
and gate_731(n997,n267,pi129);
not gate_732(n998,n997);
and gate_733(n999,n996,n998);
not gate_734(n1000,n999);
and gate_735(n1001,n266,n1000);
not gate_736(n1002,n1001);
and gate_737(n1003,n994,n1002);
not gate_738(n1004,n1003);
and gate_739(n1005,pi087,n1004);
not gate_740(n1006,n1005);
and gate_741(n1007,n991,n1006);
not gate_742(po38,n1007);
and gate_743(n1009,n267,n307);
not gate_744(n1010,n1009);
and gate_745(n1011,pi087,n1010);
not gate_746(n1012,n1011);
and gate_747(n1013,pi000,n1012);
not gate_748(n1014,n1013);
and gate_749(n1015,pi002,pi162);
and gate_750(n1016,pi000,n1015);
not gate_751(n1017,n1016);
and gate_752(n1018,pi002,pi098);
not gate_753(n1019,n1018);
and gate_754(n1020,n267,pi130);
not gate_755(n1021,n1020);
and gate_756(n1022,n1019,n1021);
not gate_757(n1023,n1022);
and gate_758(n1024,n266,n1023);
not gate_759(n1025,n1024);
and gate_760(n1026,n1017,n1025);
not gate_761(n1027,n1026);
and gate_762(n1028,pi087,n1027);
not gate_763(n1029,n1028);
and gate_764(n1030,n1014,n1029);
not gate_765(po39,n1030);
and gate_766(n1032,n267,n308);
not gate_767(n1033,n1032);
and gate_768(n1034,pi087,n1033);
not gate_769(n1035,n1034);
and gate_770(n1036,pi000,n1035);
not gate_771(n1037,n1036);
and gate_772(n1038,pi002,pi163);
and gate_773(n1039,pi000,n1038);
not gate_774(n1040,n1039);
and gate_775(n1041,pi002,pi099);
not gate_776(n1042,n1041);
and gate_777(n1043,n267,pi131);
not gate_778(n1044,n1043);
and gate_779(n1045,n1042,n1044);
not gate_780(n1046,n1045);
and gate_781(n1047,n266,n1046);
not gate_782(n1048,n1047);
and gate_783(n1049,n1040,n1048);
not gate_784(n1050,n1049);
and gate_785(n1051,pi087,n1050);
not gate_786(n1052,n1051);
and gate_787(n1053,n1037,n1052);
not gate_788(po40,n1053);
and gate_789(n1055,n267,n309);
not gate_790(n1056,n1055);
and gate_791(n1057,pi087,n1056);
not gate_792(n1058,n1057);
and gate_793(n1059,pi000,n1058);
not gate_794(n1060,n1059);
and gate_795(n1061,pi002,pi164);
and gate_796(n1062,pi000,n1061);
not gate_797(n1063,n1062);
and gate_798(n1064,pi002,pi100);
not gate_799(n1065,n1064);
and gate_800(n1066,n267,pi132);
not gate_801(n1067,n1066);
and gate_802(n1068,n1065,n1067);
not gate_803(n1069,n1068);
and gate_804(n1070,n266,n1069);
not gate_805(n1071,n1070);
and gate_806(n1072,n1063,n1071);
not gate_807(n1073,n1072);
and gate_808(n1074,pi087,n1073);
not gate_809(n1075,n1074);
and gate_810(n1076,n1060,n1075);
not gate_811(po41,n1076);
and gate_812(n1078,n267,n310);
not gate_813(n1079,n1078);
and gate_814(n1080,pi087,n1079);
not gate_815(n1081,n1080);
and gate_816(n1082,pi000,n1081);
not gate_817(n1083,n1082);
and gate_818(n1084,pi002,pi165);
and gate_819(n1085,pi000,n1084);
not gate_820(n1086,n1085);
and gate_821(n1087,pi002,pi101);
not gate_822(n1088,n1087);
and gate_823(n1089,n267,pi133);
not gate_824(n1090,n1089);
and gate_825(n1091,n1088,n1090);
not gate_826(n1092,n1091);
and gate_827(n1093,n266,n1092);
not gate_828(n1094,n1093);
and gate_829(n1095,n1086,n1094);
not gate_830(n1096,n1095);
and gate_831(n1097,pi087,n1096);
not gate_832(n1098,n1097);
and gate_833(n1099,n1083,n1098);
not gate_834(po42,n1099);
and gate_835(n1101,n267,n311);
not gate_836(n1102,n1101);
and gate_837(n1103,pi087,n1102);
not gate_838(n1104,n1103);
and gate_839(n1105,pi000,n1104);
not gate_840(n1106,n1105);
and gate_841(n1107,pi002,pi166);
and gate_842(n1108,pi000,n1107);
not gate_843(n1109,n1108);
and gate_844(n1110,pi002,pi102);
not gate_845(n1111,n1110);
and gate_846(n1112,n267,pi134);
not gate_847(n1113,n1112);
and gate_848(n1114,n1111,n1113);
not gate_849(n1115,n1114);
and gate_850(n1116,n266,n1115);
not gate_851(n1117,n1116);
and gate_852(n1118,n1109,n1117);
not gate_853(n1119,n1118);
and gate_854(n1120,pi087,n1119);
not gate_855(n1121,n1120);
and gate_856(n1122,n1106,n1121);
not gate_857(po43,n1122);
and gate_858(n1124,n267,n312);
not gate_859(n1125,n1124);
and gate_860(n1126,pi087,n1125);
not gate_861(n1127,n1126);
and gate_862(n1128,pi000,n1127);
not gate_863(n1129,n1128);
and gate_864(n1130,pi002,pi167);
and gate_865(n1131,pi000,n1130);
not gate_866(n1132,n1131);
and gate_867(n1133,pi002,pi103);
not gate_868(n1134,n1133);
and gate_869(n1135,n267,pi135);
not gate_870(n1136,n1135);
and gate_871(n1137,n1134,n1136);
not gate_872(n1138,n1137);
and gate_873(n1139,n266,n1138);
not gate_874(n1140,n1139);
and gate_875(n1141,n1132,n1140);
not gate_876(n1142,n1141);
and gate_877(n1143,pi087,n1142);
not gate_878(n1144,n1143);
and gate_879(n1145,n1129,n1144);
not gate_880(po44,n1145);
and gate_881(n1147,n267,n313);
not gate_882(n1148,n1147);
and gate_883(n1149,pi087,n1148);
not gate_884(n1150,n1149);
and gate_885(n1151,pi000,n1150);
not gate_886(n1152,n1151);
and gate_887(n1153,pi002,pi168);
and gate_888(n1154,pi000,n1153);
not gate_889(n1155,n1154);
and gate_890(n1156,pi002,pi104);
not gate_891(n1157,n1156);
and gate_892(n1158,n267,pi136);
not gate_893(n1159,n1158);
and gate_894(n1160,n1157,n1159);
not gate_895(n1161,n1160);
and gate_896(n1162,n266,n1161);
not gate_897(n1163,n1162);
and gate_898(n1164,n1155,n1163);
not gate_899(n1165,n1164);
and gate_900(n1166,pi087,n1165);
not gate_901(n1167,n1166);
and gate_902(n1168,n1152,n1167);
not gate_903(po45,n1168);
and gate_904(n1170,n267,n314);
not gate_905(n1171,n1170);
and gate_906(n1172,pi087,n1171);
not gate_907(n1173,n1172);
and gate_908(n1174,pi000,n1173);
not gate_909(n1175,n1174);
and gate_910(n1176,pi002,pi169);
and gate_911(n1177,pi000,n1176);
not gate_912(n1178,n1177);
and gate_913(n1179,pi002,pi105);
not gate_914(n1180,n1179);
and gate_915(n1181,n267,pi137);
not gate_916(n1182,n1181);
and gate_917(n1183,n1180,n1182);
not gate_918(n1184,n1183);
and gate_919(n1185,n266,n1184);
not gate_920(n1186,n1185);
and gate_921(n1187,n1178,n1186);
not gate_922(n1188,n1187);
and gate_923(n1189,pi087,n1188);
not gate_924(n1190,n1189);
and gate_925(n1191,n1175,n1190);
not gate_926(po46,n1191);
and gate_927(n1193,n267,n315);
not gate_928(n1194,n1193);
and gate_929(n1195,pi087,n1194);
not gate_930(n1196,n1195);
and gate_931(n1197,pi000,n1196);
not gate_932(n1198,n1197);
and gate_933(n1199,pi002,pi170);
and gate_934(n1200,pi000,n1199);
not gate_935(n1201,n1200);
and gate_936(n1202,pi002,pi106);
not gate_937(n1203,n1202);
and gate_938(n1204,n267,pi138);
not gate_939(n1205,n1204);
and gate_940(n1206,n1203,n1205);
not gate_941(n1207,n1206);
and gate_942(n1208,n266,n1207);
not gate_943(n1209,n1208);
and gate_944(n1210,n1201,n1209);
not gate_945(n1211,n1210);
and gate_946(n1212,pi087,n1211);
not gate_947(n1213,n1212);
and gate_948(n1214,n1198,n1213);
not gate_949(po47,n1214);
and gate_950(n1216,n267,n316);
not gate_951(n1217,n1216);
and gate_952(n1218,pi087,n1217);
not gate_953(n1219,n1218);
and gate_954(n1220,pi000,n1219);
not gate_955(n1221,n1220);
and gate_956(n1222,pi002,pi171);
and gate_957(n1223,pi000,n1222);
not gate_958(n1224,n1223);
and gate_959(n1225,pi002,pi107);
not gate_960(n1226,n1225);
and gate_961(n1227,n267,pi139);
not gate_962(n1228,n1227);
and gate_963(n1229,n1226,n1228);
not gate_964(n1230,n1229);
and gate_965(n1231,n266,n1230);
not gate_966(n1232,n1231);
and gate_967(n1233,n1224,n1232);
not gate_968(n1234,n1233);
and gate_969(n1235,pi087,n1234);
not gate_970(n1236,n1235);
and gate_971(n1237,n1221,n1236);
not gate_972(po48,n1237);
and gate_973(n1239,n267,n317);
not gate_974(n1240,n1239);
and gate_975(n1241,pi087,n1240);
not gate_976(n1242,n1241);
and gate_977(n1243,pi000,n1242);
not gate_978(n1244,n1243);
and gate_979(n1245,pi002,pi172);
and gate_980(n1246,pi000,n1245);
not gate_981(n1247,n1246);
and gate_982(n1248,pi002,pi108);
not gate_983(n1249,n1248);
and gate_984(n1250,n267,pi140);
not gate_985(n1251,n1250);
and gate_986(n1252,n1249,n1251);
not gate_987(n1253,n1252);
and gate_988(n1254,n266,n1253);
not gate_989(n1255,n1254);
and gate_990(n1256,n1247,n1255);
not gate_991(n1257,n1256);
and gate_992(n1258,pi087,n1257);
not gate_993(n1259,n1258);
and gate_994(n1260,n1244,n1259);
not gate_995(po49,n1260);
and gate_996(n1262,n267,n318);
not gate_997(n1263,n1262);
and gate_998(n1264,pi087,n1263);
not gate_999(n1265,n1264);
and gate_1000(n1266,pi000,n1265);
not gate_1001(n1267,n1266);
and gate_1002(n1268,pi002,pi173);
and gate_1003(n1269,pi000,n1268);
not gate_1004(n1270,n1269);
and gate_1005(n1271,pi002,pi109);
not gate_1006(n1272,n1271);
and gate_1007(n1273,n267,pi141);
not gate_1008(n1274,n1273);
and gate_1009(n1275,n1272,n1274);
not gate_1010(n1276,n1275);
and gate_1011(n1277,n266,n1276);
not gate_1012(n1278,n1277);
and gate_1013(n1279,n1270,n1278);
not gate_1014(n1280,n1279);
and gate_1015(n1281,pi087,n1280);
not gate_1016(n1282,n1281);
and gate_1017(n1283,n1267,n1282);
not gate_1018(po50,n1283);
and gate_1019(n1285,n267,n319);
not gate_1020(n1286,n1285);
and gate_1021(n1287,pi087,n1286);
not gate_1022(n1288,n1287);
and gate_1023(n1289,pi000,n1288);
not gate_1024(n1290,n1289);
and gate_1025(n1291,pi002,pi174);
and gate_1026(n1292,pi000,n1291);
not gate_1027(n1293,n1292);
and gate_1028(n1294,pi002,pi110);
not gate_1029(n1295,n1294);
and gate_1030(n1296,n267,pi142);
not gate_1031(n1297,n1296);
and gate_1032(n1298,n1295,n1297);
not gate_1033(n1299,n1298);
and gate_1034(n1300,n266,n1299);
not gate_1035(n1301,n1300);
and gate_1036(n1302,n1293,n1301);
not gate_1037(n1303,n1302);
and gate_1038(n1304,pi087,n1303);
not gate_1039(n1305,n1304);
and gate_1040(n1306,n1290,n1305);
not gate_1041(po51,n1306);
and gate_1042(n1308,n267,n320);
not gate_1043(n1309,n1308);
and gate_1044(n1310,pi087,n1309);
not gate_1045(n1311,n1310);
and gate_1046(n1312,pi000,n1311);
not gate_1047(n1313,n1312);
and gate_1048(n1314,pi002,pi175);
and gate_1049(n1315,pi000,n1314);
not gate_1050(n1316,n1315);
and gate_1051(n1317,pi002,pi111);
not gate_1052(n1318,n1317);
and gate_1053(n1319,n267,pi143);
not gate_1054(n1320,n1319);
and gate_1055(n1321,n1318,n1320);
not gate_1056(n1322,n1321);
and gate_1057(n1323,n266,n1322);
not gate_1058(n1324,n1323);
and gate_1059(n1325,n1316,n1324);
not gate_1060(n1326,n1325);
and gate_1061(n1327,pi087,n1326);
not gate_1062(n1328,n1327);
and gate_1063(n1329,n1313,n1328);
not gate_1064(po52,n1329);
and gate_1065(n1331,n267,n321);
not gate_1066(n1332,n1331);
and gate_1067(n1333,pi087,n1332);
not gate_1068(n1334,n1333);
and gate_1069(n1335,pi000,n1334);
not gate_1070(n1336,n1335);
and gate_1071(n1337,pi002,pi176);
and gate_1072(n1338,pi000,n1337);
not gate_1073(n1339,n1338);
and gate_1074(n1340,pi002,pi112);
not gate_1075(n1341,n1340);
and gate_1076(n1342,n267,pi144);
not gate_1077(n1343,n1342);
and gate_1078(n1344,n1341,n1343);
not gate_1079(n1345,n1344);
and gate_1080(n1346,n266,n1345);
not gate_1081(n1347,n1346);
and gate_1082(n1348,n1339,n1347);
not gate_1083(n1349,n1348);
and gate_1084(n1350,pi087,n1349);
not gate_1085(n1351,n1350);
and gate_1086(n1352,n1336,n1351);
not gate_1087(po53,n1352);
and gate_1088(n1354,n267,n322);
not gate_1089(n1355,n1354);
and gate_1090(n1356,pi087,n1355);
not gate_1091(n1357,n1356);
and gate_1092(n1358,pi000,n1357);
not gate_1093(n1359,n1358);
and gate_1094(n1360,pi002,pi177);
and gate_1095(n1361,pi000,n1360);
not gate_1096(n1362,n1361);
and gate_1097(n1363,pi002,pi113);
not gate_1098(n1364,n1363);
and gate_1099(n1365,n267,pi145);
not gate_1100(n1366,n1365);
and gate_1101(n1367,n1364,n1366);
not gate_1102(n1368,n1367);
and gate_1103(n1369,n266,n1368);
not gate_1104(n1370,n1369);
and gate_1105(n1371,n1362,n1370);
not gate_1106(n1372,n1371);
and gate_1107(n1373,pi087,n1372);
not gate_1108(n1374,n1373);
and gate_1109(n1375,n1359,n1374);
not gate_1110(po54,n1375);
and gate_1111(n1377,n267,n323);
not gate_1112(n1378,n1377);
and gate_1113(n1379,pi087,n1378);
not gate_1114(n1380,n1379);
and gate_1115(n1381,pi000,n1380);
not gate_1116(n1382,n1381);
and gate_1117(n1383,pi002,pi178);
and gate_1118(n1384,pi000,n1383);
not gate_1119(n1385,n1384);
and gate_1120(n1386,pi002,pi114);
not gate_1121(n1387,n1386);
and gate_1122(n1388,n267,pi146);
not gate_1123(n1389,n1388);
and gate_1124(n1390,n1387,n1389);
not gate_1125(n1391,n1390);
and gate_1126(n1392,n266,n1391);
not gate_1127(n1393,n1392);
and gate_1128(n1394,n1385,n1393);
not gate_1129(n1395,n1394);
and gate_1130(n1396,pi087,n1395);
not gate_1131(n1397,n1396);
and gate_1132(n1398,n1382,n1397);
not gate_1133(po55,n1398);
and gate_1134(n1400,n267,n324);
not gate_1135(n1401,n1400);
and gate_1136(n1402,pi087,n1401);
not gate_1137(n1403,n1402);
and gate_1138(n1404,pi000,n1403);
not gate_1139(n1405,n1404);
and gate_1140(n1406,pi002,pi179);
and gate_1141(n1407,pi000,n1406);
not gate_1142(n1408,n1407);
and gate_1143(n1409,pi002,pi115);
not gate_1144(n1410,n1409);
and gate_1145(n1411,n267,pi147);
not gate_1146(n1412,n1411);
and gate_1147(n1413,n1410,n1412);
not gate_1148(n1414,n1413);
and gate_1149(n1415,n266,n1414);
not gate_1150(n1416,n1415);
and gate_1151(n1417,n1408,n1416);
not gate_1152(n1418,n1417);
and gate_1153(n1419,pi087,n1418);
not gate_1154(n1420,n1419);
and gate_1155(n1421,n1405,n1420);
not gate_1156(po56,n1421);
and gate_1157(n1423,n267,n325);
not gate_1158(n1424,n1423);
and gate_1159(n1425,pi087,n1424);
not gate_1160(n1426,n1425);
and gate_1161(n1427,pi000,n1426);
not gate_1162(n1428,n1427);
and gate_1163(n1429,pi002,pi180);
and gate_1164(n1430,pi000,n1429);
not gate_1165(n1431,n1430);
and gate_1166(n1432,pi002,pi116);
not gate_1167(n1433,n1432);
and gate_1168(n1434,n267,pi148);
not gate_1169(n1435,n1434);
and gate_1170(n1436,n1433,n1435);
not gate_1171(n1437,n1436);
and gate_1172(n1438,n266,n1437);
not gate_1173(n1439,n1438);
and gate_1174(n1440,n1431,n1439);
not gate_1175(n1441,n1440);
and gate_1176(n1442,pi087,n1441);
not gate_1177(n1443,n1442);
and gate_1178(n1444,n1428,n1443);
not gate_1179(po57,n1444);
and gate_1180(n1446,n267,n326);
not gate_1181(n1447,n1446);
and gate_1182(n1448,pi087,n1447);
not gate_1183(n1449,n1448);
and gate_1184(n1450,pi000,n1449);
not gate_1185(n1451,n1450);
and gate_1186(n1452,pi002,pi181);
and gate_1187(n1453,pi000,n1452);
not gate_1188(n1454,n1453);
and gate_1189(n1455,pi002,pi117);
not gate_1190(n1456,n1455);
and gate_1191(n1457,n267,pi149);
not gate_1192(n1458,n1457);
and gate_1193(n1459,n1456,n1458);
not gate_1194(n1460,n1459);
and gate_1195(n1461,n266,n1460);
not gate_1196(n1462,n1461);
and gate_1197(n1463,n1454,n1462);
not gate_1198(n1464,n1463);
and gate_1199(n1465,pi087,n1464);
not gate_1200(n1466,n1465);
and gate_1201(n1467,n1451,n1466);
not gate_1202(po58,n1467);
and gate_1203(n1469,n267,n327);
not gate_1204(n1470,n1469);
and gate_1205(n1471,pi087,n1470);
not gate_1206(n1472,n1471);
and gate_1207(n1473,pi000,n1472);
not gate_1208(n1474,n1473);
and gate_1209(n1475,pi002,pi182);
and gate_1210(n1476,pi000,n1475);
not gate_1211(n1477,n1476);
and gate_1212(n1478,pi002,pi118);
not gate_1213(n1479,n1478);
and gate_1214(n1480,n267,pi150);
not gate_1215(n1481,n1480);
and gate_1216(n1482,n1479,n1481);
not gate_1217(n1483,n1482);
and gate_1218(n1484,n266,n1483);
not gate_1219(n1485,n1484);
and gate_1220(n1486,n1477,n1485);
not gate_1221(n1487,n1486);
and gate_1222(n1488,pi087,n1487);
not gate_1223(n1489,n1488);
and gate_1224(n1490,n1474,n1489);
not gate_1225(po59,n1490);
and gate_1226(n1492,pi184,pi188);
and gate_1227(po60,n267,n1492);
and gate_1228(n1494,pi000,n328);
not gate_1229(n1495,n1494);
and gate_1230(n1496,n267,pi189);
not gate_1231(n1497,n1496);
and gate_1232(n1498,n266,n1496);
and gate_1233(n1499,pi184,n1498);
not gate_1234(n1500,n1499);
and gate_1235(n1501,n1495,n1500);
and gate_1236(n1502,pi000,pi184);
and gate_1237(n1503,n1497,n1502);
not gate_1238(n1504,n1503);
and gate_1239(n1505,n1501,n1504);
not gate_1240(po61,n1505);
and gate_1241(n1507,n267,pi190);
not gate_1242(n1508,n1507);
and gate_1243(n1509,n266,n1507);
and gate_1244(n1510,pi184,n1509);
not gate_1245(n1511,n1510);
and gate_1246(n1512,n1495,n1511);
and gate_1247(n1513,n1502,n1508);
not gate_1248(n1514,n1513);
and gate_1249(n1515,n1512,n1514);
not gate_1250(po62,n1515);
and gate_1251(n1517,n267,n332);
and gate_1252(n1518,n1502,n1517);
not gate_1253(n1519,n1518);
and gate_1254(n1520,n1495,n1519);
and gate_1255(n1521,pi002,n1502);
and gate_1256(n1522,pi195,n1521);
not gate_1257(n1523,n1522);
and gate_1258(n1524,n266,pi184);
and gate_1259(n1525,pi002,pi183);
not gate_1260(n1526,n1525);
and gate_1261(n1527,n267,pi191);
not gate_1262(n1528,n1527);
and gate_1263(n1529,n1526,n1528);
not gate_1264(n1530,n1529);
and gate_1265(n1531,n1524,n1530);
not gate_1266(n1532,n1531);
and gate_1267(n1533,n1523,n1532);
and gate_1268(n1534,n1520,n1533);
not gate_1269(po63,n1534);
and gate_1270(n1536,n267,n333);
not gate_1271(n1537,n1536);
and gate_1272(n1538,n1502,n1536);
not gate_1273(n1539,n1538);
and gate_1274(n1540,n1495,n1539);
and gate_1275(n1541,pi196,n1521);
not gate_1276(n1542,n1541);
and gate_1277(n1543,n1524,n1537);
and gate_1278(n1544,pi002,n329);
not gate_1279(n1545,n1544);
and gate_1280(n1546,n1543,n1545);
not gate_1281(n1547,n1546);
and gate_1282(n1548,n1542,n1547);
and gate_1283(n1549,n1540,n1548);
not gate_1284(po64,n1549);
and gate_1285(n1551,n267,n334);
not gate_1286(n1552,n1551);
and gate_1287(n1553,n1502,n1551);
not gate_1288(n1554,n1553);
and gate_1289(n1555,n1495,n1554);
and gate_1290(n1556,pi197,n1521);
not gate_1291(n1557,n1556);
and gate_1292(n1558,n1524,n1552);
and gate_1293(n1559,pi002,n330);
not gate_1294(n1560,n1559);
and gate_1295(n1561,n1558,n1560);
not gate_1296(n1562,n1561);
and gate_1297(n1563,n1557,n1562);
and gate_1298(n1564,n1555,n1563);
not gate_1299(po65,n1564);
and gate_1300(n1566,n267,n335);
not gate_1301(n1567,n1566);
and gate_1302(n1568,n1502,n1566);
not gate_1303(n1569,n1568);
and gate_1304(n1570,n1495,n1569);
and gate_1305(n1571,pi198,n1521);
not gate_1306(n1572,n1571);
and gate_1307(n1573,n1524,n1567);
and gate_1308(n1574,pi002,n331);
not gate_1309(n1575,n1574);
and gate_1310(n1576,n1573,n1575);
not gate_1311(n1577,n1576);
and gate_1312(n1578,n1572,n1577);
and gate_1313(n1579,n1570,n1578);
not gate_1314(po66,n1579);
endmodule
