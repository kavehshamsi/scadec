
module c432_xrnd_8 ( G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, 
        G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, 
        G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, 
        G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, 
        G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, 
        G431gat, G432gat, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7 );
  input G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat,
         G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat,
         G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat,
         G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat,
         G108gat, G112gat, G115gat, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7;
  output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
  wire   n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270;

  NAND2_X1 U144 ( .A1(n143), .A2(n144), .ZN(G432gat) );
  NAND2_X1 U145 ( .A1(n145), .A2(n146), .ZN(n144) );
  NAND3_X1 U146 ( .A1(n147), .A2(n148), .A3(n149), .ZN(n145) );
  NAND3_X1 U147 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n147) );
  NAND4_X1 U148 ( .A1(n153), .A2(n143), .A3(n146), .A4(n148), .ZN(G431gat) );
  NAND2_X1 U149 ( .A1(n154), .A2(n155), .ZN(n148) );
  INV_X1 U150 ( .A(n156), .ZN(n154) );
  OR2_X1 U151 ( .A1(n151), .A2(n156), .ZN(n153) );
  NAND4_X1 U152 ( .A1(n149), .A2(n157), .A3(n143), .A4(n146), .ZN(G430gat) );
  XOR2_X1 U153 ( .A(n150), .B(keyinput7), .Z(n149) );
  NOR2_X1 U154 ( .A1(n158), .A2(n159), .ZN(G421gat) );
  NOR4_X1 U155 ( .A1(n160), .A2(n161), .A3(n162), .A4(n163), .ZN(n159) );
  AND2_X1 U156 ( .A1(G370gat), .A2(G14gat), .ZN(n162) );
  AND2_X1 U157 ( .A1(G329gat), .A2(G8gat), .ZN(n161) );
  NOR2_X1 U158 ( .A1(n164), .A2(n165), .ZN(n160) );
  NOR4_X1 U159 ( .A1(n166), .A2(n152), .A3(n155), .A4(n156), .ZN(n158) );
  NAND2_X1 U160 ( .A1(n157), .A2(n150), .ZN(n156) );
  NAND3_X1 U161 ( .A1(n167), .A2(n168), .A3(n169), .ZN(n150) );
  NAND2_X1 U162 ( .A1(G53gat), .A2(G370gat), .ZN(n169) );
  NAND2_X1 U163 ( .A1(n170), .A2(n171), .ZN(n168) );
  NAND2_X1 U164 ( .A1(G43gat), .A2(n164), .ZN(n170) );
  NAND2_X1 U165 ( .A1(G47gat), .A2(G329gat), .ZN(n167) );
  NAND3_X1 U166 ( .A1(n172), .A2(n173), .A3(n174), .ZN(n157) );
  NAND2_X1 U167 ( .A1(G60gat), .A2(G329gat), .ZN(n173) );
  NAND2_X1 U168 ( .A1(G66gat), .A2(G370gat), .ZN(n172) );
  AND3_X1 U169 ( .A1(n175), .A2(n176), .A3(n177), .ZN(n155) );
  NAND2_X1 U170 ( .A1(G73gat), .A2(G329gat), .ZN(n176) );
  NAND2_X1 U171 ( .A1(G79gat), .A2(G370gat), .ZN(n175) );
  XNOR2_X1 U172 ( .A(n178), .B(keyinput5), .ZN(n152) );
  NAND4_X1 U173 ( .A1(G95gat), .A2(n179), .A3(n180), .A4(n181), .ZN(n178) );
  NAND2_X1 U174 ( .A1(G99gat), .A2(G329gat), .ZN(n180) );
  NAND2_X1 U175 ( .A1(G105gat), .A2(G370gat), .ZN(n179) );
  NAND4_X1 U176 ( .A1(n151), .A2(n143), .A3(n146), .A4(n182), .ZN(n166) );
  NAND4_X1 U177 ( .A1(G108gat), .A2(n183), .A3(n184), .A4(n185), .ZN(n182) );
  NAND2_X1 U178 ( .A1(G115gat), .A2(G370gat), .ZN(n184) );
  NAND4_X1 U179 ( .A1(n186), .A2(G30gat), .A3(n187), .A4(n188), .ZN(n146) );
  NAND2_X1 U180 ( .A1(G34gat), .A2(G329gat), .ZN(n188) );
  NAND2_X1 U181 ( .A1(G40gat), .A2(G370gat), .ZN(n187) );
  MUX2_X1 U182 ( .A(n189), .B(n190), .S(keyinput6), .Z(n186) );
  NOR2_X1 U183 ( .A1(n164), .A2(n191), .ZN(n190) );
  INV_X1 U184 ( .A(G223gat), .ZN(n164) );
  NAND4_X1 U185 ( .A1(G17gat), .A2(n192), .A3(n193), .A4(n194), .ZN(n143) );
  NAND2_X1 U186 ( .A1(G21gat), .A2(G329gat), .ZN(n193) );
  NAND2_X1 U187 ( .A1(G27gat), .A2(G370gat), .ZN(n192) );
  NAND4_X1 U188 ( .A1(G82gat), .A2(n195), .A3(n196), .A4(n197), .ZN(n151) );
  OR2_X1 U189 ( .A1(n198), .A2(n199), .ZN(n196) );
  NAND2_X1 U190 ( .A1(G92gat), .A2(G370gat), .ZN(n195) );
  NAND4_X1 U191 ( .A1(n200), .A2(n201), .A3(n202), .A4(n203), .ZN(G370gat) );
  NOR3_X1 U192 ( .A1(n204), .A2(n205), .A3(n206), .ZN(n203) );
  NOR3_X1 U193 ( .A1(n207), .A2(G40gat), .A3(G34gat), .ZN(n206) );
  NOR3_X1 U194 ( .A1(n208), .A2(G27gat), .A3(G21gat), .ZN(n205) );
  NAND3_X1 U195 ( .A1(n209), .A2(n210), .A3(n211), .ZN(n204) );
  NAND4_X1 U196 ( .A1(G108gat), .A2(n183), .A3(n185), .A4(n212), .ZN(n211) );
  INV_X1 U197 ( .A(G115gat), .ZN(n212) );
  NAND2_X1 U198 ( .A1(G112gat), .A2(G329gat), .ZN(n185) );
  NAND3_X1 U199 ( .A1(n213), .A2(n214), .A3(n177), .ZN(n210) );
  INV_X1 U200 ( .A(n215), .ZN(n177) );
  INV_X1 U201 ( .A(G79gat), .ZN(n214) );
  NAND2_X1 U202 ( .A1(G329gat), .A2(n216), .ZN(n213) );
  NAND3_X1 U203 ( .A1(n217), .A2(n218), .A3(n174), .ZN(n209) );
  INV_X1 U204 ( .A(n219), .ZN(n174) );
  INV_X1 U205 ( .A(G66gat), .ZN(n218) );
  NAND2_X1 U206 ( .A1(G329gat), .A2(n220), .ZN(n217) );
  NOR3_X1 U207 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n202) );
  NOR3_X1 U208 ( .A1(n224), .A2(G8gat), .A3(G14gat), .ZN(n223) );
  NOR3_X1 U209 ( .A1(n225), .A2(G53gat), .A3(G47gat), .ZN(n222) );
  NOR3_X1 U210 ( .A1(n226), .A2(G99gat), .A3(G105gat), .ZN(n221) );
  NAND2_X1 U211 ( .A1(n227), .A2(n199), .ZN(n201) );
  INV_X1 U212 ( .A(G329gat), .ZN(n199) );
  NAND3_X1 U213 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n227) );
  NOR3_X1 U214 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n230) );
  NOR2_X1 U215 ( .A1(G40gat), .A2(n207), .ZN(n233) );
  NOR2_X1 U216 ( .A1(G27gat), .A2(n208), .ZN(n232) );
  NOR2_X1 U217 ( .A1(G53gat), .A2(n225), .ZN(n231) );
  OR2_X1 U218 ( .A1(n224), .A2(G14gat), .ZN(n229) );
  OR2_X1 U219 ( .A1(n226), .A2(G105gat), .ZN(n228) );
  XOR2_X1 U220 ( .A(n234), .B(keyinput0), .Z(n200) );
  NAND4_X1 U221 ( .A1(G82gat), .A2(n235), .A3(n197), .A4(n236), .ZN(n234) );
  INV_X1 U222 ( .A(G92gat), .ZN(n236) );
  NAND2_X1 U223 ( .A1(G329gat), .A2(n237), .ZN(n235) );
  NAND4_X1 U224 ( .A1(n238), .A2(n239), .A3(n240), .A4(n241), .ZN(G329gat) );
  NOR4_X1 U225 ( .A1(n242), .A2(n243), .A3(n244), .A4(n245), .ZN(n241) );
  NOR2_X1 U226 ( .A1(G99gat), .A2(n226), .ZN(n245) );
  NAND2_X1 U227 ( .A1(G95gat), .A2(n181), .ZN(n226) );
  NAND2_X1 U228 ( .A1(G223gat), .A2(n246), .ZN(n181) );
  NOR2_X1 U229 ( .A1(G8gat), .A2(n224), .ZN(n244) );
  NAND2_X1 U230 ( .A1(n247), .A2(n248), .ZN(n224) );
  NAND2_X1 U231 ( .A1(G223gat), .A2(n249), .ZN(n248) );
  NAND2_X1 U232 ( .A1(G4gat), .A2(n165), .ZN(n249) );
  INV_X1 U233 ( .A(G1gat), .ZN(n165) );
  XOR2_X1 U234 ( .A(keyinput3), .B(G4gat), .Z(n247) );
  NOR2_X1 U235 ( .A1(G47gat), .A2(n225), .ZN(n243) );
  NAND2_X1 U236 ( .A1(G43gat), .A2(n250), .ZN(n225) );
  XOR2_X1 U237 ( .A(G223gat), .B(n251), .Z(n250) );
  XOR2_X1 U238 ( .A(n171), .B(keyinput2), .Z(n251) );
  NOR2_X1 U239 ( .A1(G34gat), .A2(n207), .ZN(n242) );
  NAND2_X1 U240 ( .A1(G30gat), .A2(n189), .ZN(n207) );
  NAND2_X1 U241 ( .A1(G223gat), .A2(n252), .ZN(n189) );
  AND3_X1 U242 ( .A1(n216), .A2(n237), .A3(n220), .ZN(n240) );
  OR2_X1 U243 ( .A1(n219), .A2(G60gat), .ZN(n220) );
  NAND2_X1 U244 ( .A1(G56gat), .A2(n253), .ZN(n219) );
  NAND2_X1 U245 ( .A1(G50gat), .A2(G223gat), .ZN(n253) );
  NAND3_X1 U246 ( .A1(G82gat), .A2(n197), .A3(n198), .ZN(n237) );
  XNOR2_X1 U247 ( .A(keyinput4), .B(G86gat), .ZN(n198) );
  NAND2_X1 U248 ( .A1(G223gat), .A2(n254), .ZN(n197) );
  OR2_X1 U249 ( .A1(n215), .A2(G73gat), .ZN(n216) );
  NAND2_X1 U250 ( .A1(G69gat), .A2(n255), .ZN(n215) );
  NAND2_X1 U251 ( .A1(G63gat), .A2(G223gat), .ZN(n255) );
  NAND3_X1 U252 ( .A1(n183), .A2(n256), .A3(G108gat), .ZN(n239) );
  INV_X1 U253 ( .A(G112gat), .ZN(n256) );
  NAND2_X1 U254 ( .A1(G102gat), .A2(G223gat), .ZN(n183) );
  OR2_X1 U255 ( .A1(n208), .A2(G21gat), .ZN(n238) );
  NAND2_X1 U256 ( .A1(G17gat), .A2(n194), .ZN(n208) );
  NAND2_X1 U257 ( .A1(G11gat), .A2(G223gat), .ZN(n194) );
  NAND4_X1 U258 ( .A1(n257), .A2(n254), .A3(n258), .A4(n259), .ZN(G223gat) );
  NOR4_X1 U259 ( .A1(n260), .A2(n261), .A3(n262), .A4(n263), .ZN(n259) );
  NOR2_X1 U260 ( .A1(G63gat), .A2(n264), .ZN(n263) );
  INV_X1 U261 ( .A(G69gat), .ZN(n264) );
  NOR2_X1 U262 ( .A1(G50gat), .A2(n265), .ZN(n262) );
  INV_X1 U263 ( .A(G56gat), .ZN(n265) );
  NOR2_X1 U264 ( .A1(G1gat), .A2(n163), .ZN(n261) );
  INV_X1 U265 ( .A(G4gat), .ZN(n163) );
  NOR2_X1 U266 ( .A1(G11gat), .A2(n266), .ZN(n260) );
  INV_X1 U267 ( .A(G17gat), .ZN(n266) );
  AND3_X1 U268 ( .A1(n246), .A2(n171), .A3(n252), .ZN(n258) );
  NAND2_X1 U269 ( .A1(G30gat), .A2(n191), .ZN(n252) );
  INV_X1 U270 ( .A(G24gat), .ZN(n191) );
  NAND2_X1 U271 ( .A1(n267), .A2(G43gat), .ZN(n171) );
  INV_X1 U272 ( .A(G37gat), .ZN(n267) );
  NAND2_X1 U273 ( .A1(n268), .A2(G95gat), .ZN(n246) );
  INV_X1 U274 ( .A(G89gat), .ZN(n268) );
  NAND2_X1 U275 ( .A1(n269), .A2(G82gat), .ZN(n254) );
  XNOR2_X1 U276 ( .A(keyinput1), .B(G76gat), .ZN(n269) );
  NAND2_X1 U277 ( .A1(G108gat), .A2(n270), .ZN(n257) );
  INV_X1 U278 ( .A(G102gat), .ZN(n270) );
endmodule

