
module c432_xrnd_16 ( G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, 
        G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, 
        G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, 
        G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, 
        G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, 
        G431gat, G432gat, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15
 );
  input G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat,
         G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat,
         G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat,
         G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat,
         G108gat, G112gat, G115gat, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15;
  output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
  wire   n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289;

  NAND2_X1 U147 ( .A1(n146), .A2(n147), .ZN(G432gat) );
  NAND2_X1 U148 ( .A1(n148), .A2(n149), .ZN(n147) );
  NAND3_X1 U149 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n148) );
  NAND2_X1 U150 ( .A1(n153), .A2(n154), .ZN(n152) );
  INV_X1 U151 ( .A(n155), .ZN(n153) );
  NAND4_X1 U152 ( .A1(n156), .A2(n157), .A3(n158), .A4(n159), .ZN(n150) );
  NAND3_X1 U153 ( .A1(n160), .A2(n149), .A3(n146), .ZN(G431gat) );
  NAND3_X1 U154 ( .A1(n151), .A2(n154), .A3(n161), .ZN(n160) );
  NOR2_X1 U155 ( .A1(n162), .A2(n163), .ZN(G421gat) );
  NOR4_X1 U156 ( .A1(G430gat), .A2(n164), .A3(n165), .A4(n161), .ZN(n163) );
  NAND2_X1 U157 ( .A1(n155), .A2(n159), .ZN(n161) );
  NAND4_X1 U158 ( .A1(G82gat), .A2(n166), .A3(n167), .A4(n168), .ZN(n159) );
  NAND2_X1 U159 ( .A1(n169), .A2(n170), .ZN(n168) );
  NAND2_X1 U160 ( .A1(G76gat), .A2(G223gat), .ZN(n167) );
  NAND2_X1 U161 ( .A1(G86gat), .A2(G329gat), .ZN(n166) );
  NAND3_X1 U162 ( .A1(n171), .A2(n172), .A3(n173), .ZN(n155) );
  NAND2_X1 U163 ( .A1(G79gat), .A2(n169), .ZN(n172) );
  NAND2_X1 U164 ( .A1(G73gat), .A2(G329gat), .ZN(n171) );
  AND3_X1 U165 ( .A1(n156), .A2(n158), .A3(n157), .ZN(n165) );
  NAND2_X1 U166 ( .A1(G99gat), .A2(G329gat), .ZN(n157) );
  NAND2_X1 U167 ( .A1(G105gat), .A2(n169), .ZN(n158) );
  AND2_X1 U168 ( .A1(G95gat), .A2(n174), .ZN(n156) );
  NOR4_X1 U169 ( .A1(n175), .A2(n176), .A3(n177), .A4(n178), .ZN(n164) );
  NOR2_X1 U170 ( .A1(n179), .A2(n180), .ZN(n176) );
  AND2_X1 U171 ( .A1(G329gat), .A2(G112gat), .ZN(n175) );
  NAND4_X1 U172 ( .A1(n146), .A2(n151), .A3(n154), .A4(n149), .ZN(G430gat) );
  NAND4_X1 U173 ( .A1(G30gat), .A2(n181), .A3(n182), .A4(n183), .ZN(n149) );
  NAND2_X1 U174 ( .A1(G40gat), .A2(n169), .ZN(n182) );
  NAND2_X1 U175 ( .A1(G34gat), .A2(G329gat), .ZN(n181) );
  NAND3_X1 U176 ( .A1(n184), .A2(n185), .A3(n186), .ZN(n154) );
  NAND2_X1 U177 ( .A1(G60gat), .A2(G329gat), .ZN(n186) );
  NAND2_X1 U178 ( .A1(n187), .A2(n188), .ZN(n185) );
  NAND2_X1 U179 ( .A1(G56gat), .A2(n189), .ZN(n187) );
  NAND2_X1 U180 ( .A1(G66gat), .A2(n169), .ZN(n184) );
  NAND4_X1 U181 ( .A1(G43gat), .A2(n190), .A3(n191), .A4(n192), .ZN(n151) );
  NAND2_X1 U182 ( .A1(n193), .A2(G329gat), .ZN(n191) );
  NAND2_X1 U183 ( .A1(G53gat), .A2(n169), .ZN(n190) );
  XOR2_X1 U184 ( .A(n194), .B(keyinput7), .Z(n146) );
  NAND4_X1 U185 ( .A1(G17gat), .A2(n195), .A3(n196), .A4(n197), .ZN(n194) );
  NAND2_X1 U186 ( .A1(G27gat), .A2(n169), .ZN(n196) );
  INV_X1 U187 ( .A(n180), .ZN(n169) );
  NAND2_X1 U188 ( .A1(G21gat), .A2(G329gat), .ZN(n195) );
  NOR4_X1 U189 ( .A1(n198), .A2(n199), .A3(n200), .A4(n201), .ZN(n162) );
  XOR2_X1 U190 ( .A(keyinput6), .B(n202), .Z(n201) );
  AND2_X1 U191 ( .A1(G223gat), .A2(G1gat), .ZN(n202) );
  NOR2_X1 U192 ( .A1(n180), .A2(n203), .ZN(n199) );
  XNOR2_X1 U193 ( .A(G370gat), .B(keyinput15), .ZN(n180) );
  AND2_X1 U194 ( .A1(G329gat), .A2(n204), .ZN(n198) );
  NAND4_X1 U195 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(G370gat) );
  NAND3_X1 U196 ( .A1(n209), .A2(n210), .A3(n173), .ZN(n208) );
  INV_X1 U197 ( .A(n211), .ZN(n173) );
  INV_X1 U198 ( .A(G79gat), .ZN(n210) );
  XNOR2_X1 U199 ( .A(n212), .B(n213), .ZN(n209) );
  NAND3_X1 U200 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n207) );
  INV_X1 U201 ( .A(G66gat), .ZN(n215) );
  XNOR2_X1 U202 ( .A(n217), .B(n218), .ZN(n214) );
  XNOR2_X1 U203 ( .A(n219), .B(keyinput0), .ZN(n218) );
  NAND4_X1 U204 ( .A1(G43gat), .A2(n220), .A3(n192), .A4(n221), .ZN(n206) );
  INV_X1 U205 ( .A(G53gat), .ZN(n221) );
  XNOR2_X1 U206 ( .A(n222), .B(n213), .ZN(n220) );
  MUX2_X1 U207 ( .A(n223), .B(n224), .S(n213), .Z(n205) );
  INV_X1 U208 ( .A(n217), .ZN(n213) );
  XNOR2_X1 U209 ( .A(G329gat), .B(keyinput4), .ZN(n217) );
  NOR4_X1 U210 ( .A1(n225), .A2(n226), .A3(n227), .A4(n228), .ZN(n224) );
  NOR2_X1 U211 ( .A1(G105gat), .A2(n229), .ZN(n228) );
  AND2_X1 U212 ( .A1(n203), .A2(n230), .ZN(n227) );
  INV_X1 U213 ( .A(G14gat), .ZN(n203) );
  NOR2_X1 U214 ( .A1(n231), .A2(n232), .ZN(n226) );
  INV_X1 U215 ( .A(n233), .ZN(n232) );
  NAND3_X1 U216 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n225) );
  NAND2_X1 U217 ( .A1(n237), .A2(n179), .ZN(n236) );
  OR2_X1 U218 ( .A1(n238), .A2(n170), .ZN(n235) );
  NAND2_X1 U219 ( .A1(n239), .A2(n240), .ZN(n234) );
  INV_X1 U220 ( .A(G27gat), .ZN(n240) );
  NOR4_X1 U221 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n223) );
  NOR3_X1 U222 ( .A1(n245), .A2(G105gat), .A3(n246), .ZN(n244) );
  NOR3_X1 U223 ( .A1(n247), .A2(G14gat), .A3(n230), .ZN(n243) );
  NOR2_X1 U224 ( .A1(n233), .A2(n231), .ZN(n242) );
  XOR2_X1 U225 ( .A(n248), .B(keyinput5), .Z(n231) );
  OR3_X1 U226 ( .A1(n249), .A2(G40gat), .A3(n250), .ZN(n248) );
  NAND3_X1 U227 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n241) );
  NAND3_X1 U228 ( .A1(n254), .A2(n255), .A3(n179), .ZN(n253) );
  XNOR2_X1 U229 ( .A(keyinput14), .B(G115gat), .ZN(n179) );
  INV_X1 U230 ( .A(n237), .ZN(n255) );
  OR3_X1 U231 ( .A1(n256), .A2(n257), .A3(n170), .ZN(n252) );
  XOR2_X1 U232 ( .A(keyinput2), .B(G92gat), .Z(n170) );
  OR3_X1 U233 ( .A1(n239), .A2(G27gat), .A3(n258), .ZN(n251) );
  NAND4_X1 U234 ( .A1(n229), .A2(n238), .A3(n259), .A4(n260), .ZN(G329gat) );
  NOR4_X1 U235 ( .A1(n237), .A2(n212), .A3(n222), .A4(n219), .ZN(n260) );
  XNOR2_X1 U236 ( .A(n261), .B(keyinput3), .ZN(n219) );
  NAND2_X1 U237 ( .A1(n216), .A2(n262), .ZN(n261) );
  INV_X1 U238 ( .A(G60gat), .ZN(n262) );
  AND2_X1 U239 ( .A1(G56gat), .A2(n263), .ZN(n216) );
  OR2_X1 U240 ( .A1(n264), .A2(n189), .ZN(n263) );
  INV_X1 U241 ( .A(G223gat), .ZN(n189) );
  AND3_X1 U242 ( .A1(n265), .A2(n192), .A3(n266), .ZN(n222) );
  XOR2_X1 U243 ( .A(keyinput9), .B(n267), .Z(n266) );
  NOR2_X1 U244 ( .A1(n268), .A2(n193), .ZN(n267) );
  XOR2_X1 U245 ( .A(keyinput11), .B(G47gat), .Z(n193) );
  NAND2_X1 U246 ( .A1(G37gat), .A2(G223gat), .ZN(n192) );
  NAND2_X1 U247 ( .A1(G223gat), .A2(n268), .ZN(n265) );
  NOR2_X1 U248 ( .A1(n211), .A2(G73gat), .ZN(n212) );
  NAND2_X1 U249 ( .A1(n269), .A2(n270), .ZN(n211) );
  NAND2_X1 U250 ( .A1(G63gat), .A2(G223gat), .ZN(n270) );
  NOR2_X1 U251 ( .A1(n271), .A2(G112gat), .ZN(n237) );
  INV_X1 U252 ( .A(n254), .ZN(n271) );
  NOR2_X1 U253 ( .A1(n178), .A2(n177), .ZN(n254) );
  AND2_X1 U254 ( .A1(G102gat), .A2(G223gat), .ZN(n177) );
  NOR3_X1 U255 ( .A1(n239), .A2(n233), .A3(n230), .ZN(n259) );
  NOR2_X1 U256 ( .A1(n247), .A2(n204), .ZN(n230) );
  XOR2_X1 U257 ( .A(keyinput10), .B(G8gat), .Z(n204) );
  NAND2_X1 U258 ( .A1(G4gat), .A2(n272), .ZN(n247) );
  NAND2_X1 U259 ( .A1(G1gat), .A2(G223gat), .ZN(n272) );
  NOR3_X1 U260 ( .A1(n249), .A2(G34gat), .A3(n250), .ZN(n233) );
  INV_X1 U261 ( .A(n183), .ZN(n249) );
  NAND2_X1 U262 ( .A1(G223gat), .A2(n273), .ZN(n183) );
  NOR2_X1 U263 ( .A1(n258), .A2(G21gat), .ZN(n239) );
  NAND2_X1 U264 ( .A1(G17gat), .A2(n197), .ZN(n258) );
  NAND2_X1 U265 ( .A1(G223gat), .A2(n274), .ZN(n197) );
  INV_X1 U266 ( .A(n257), .ZN(n238) );
  NOR2_X1 U267 ( .A1(n256), .A2(G86gat), .ZN(n257) );
  NAND2_X1 U268 ( .A1(G82gat), .A2(n275), .ZN(n256) );
  NAND2_X1 U269 ( .A1(G223gat), .A2(n276), .ZN(n275) );
  INV_X1 U270 ( .A(n246), .ZN(n229) );
  NOR2_X1 U271 ( .A1(n245), .A2(G99gat), .ZN(n246) );
  NAND2_X1 U272 ( .A1(G95gat), .A2(n174), .ZN(n245) );
  NAND2_X1 U273 ( .A1(G89gat), .A2(G223gat), .ZN(n174) );
  NAND4_X1 U274 ( .A1(n277), .A2(n278), .A3(n279), .A4(n280), .ZN(G223gat) );
  NOR4_X1 U275 ( .A1(n281), .A2(n282), .A3(n283), .A4(n264), .ZN(n280) );
  XOR2_X1 U276 ( .A(n284), .B(n188), .Z(n264) );
  NAND2_X1 U277 ( .A1(n285), .A2(G56gat), .ZN(n188) );
  INV_X1 U278 ( .A(G50gat), .ZN(n285) );
  XNOR2_X1 U279 ( .A(keyinput8), .B(keyinput13), .ZN(n284) );
  NOR2_X1 U280 ( .A1(G89gat), .A2(n286), .ZN(n283) );
  INV_X1 U281 ( .A(G95gat), .ZN(n286) );
  NOR2_X1 U282 ( .A1(G37gat), .A2(n268), .ZN(n282) );
  INV_X1 U283 ( .A(G43gat), .ZN(n268) );
  NOR2_X1 U284 ( .A1(G1gat), .A2(n200), .ZN(n281) );
  INV_X1 U285 ( .A(G4gat), .ZN(n200) );
  AND3_X1 U286 ( .A1(n276), .A2(n274), .A3(n273), .ZN(n279) );
  OR2_X1 U287 ( .A1(G24gat), .A2(n250), .ZN(n273) );
  INV_X1 U288 ( .A(G30gat), .ZN(n250) );
  NAND2_X1 U289 ( .A1(n287), .A2(G17gat), .ZN(n274) );
  INV_X1 U290 ( .A(G11gat), .ZN(n287) );
  NAND2_X1 U291 ( .A1(n288), .A2(G82gat), .ZN(n276) );
  XNOR2_X1 U292 ( .A(G76gat), .B(keyinput1), .ZN(n288) );
  NAND2_X1 U293 ( .A1(n269), .A2(n289), .ZN(n278) );
  INV_X1 U294 ( .A(G63gat), .ZN(n289) );
  XOR2_X1 U295 ( .A(keyinput12), .B(G69gat), .Z(n269) );
  OR2_X1 U296 ( .A1(n178), .A2(G102gat), .ZN(n277) );
  INV_X1 U297 ( .A(G108gat), .ZN(n178) );
endmodule

