// Verilog File 
module seq (pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
pi39,pi40,po00,po01,po02,po03,po04,po05,po06,po07,
po08,po09,po10,po11,po12,po13,po14,po15,po16,po17,
po18,po19,po20,po21,po22,po23,po24,po25,po26,po27,
po28,po29,po30,po31,po32,po33,po34);

input pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
pi39,pi40;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18,
po19,po20,po21,po22,po23,po24,po25,po26,po27,po28,
po29,po30,po31,po32,po33,po34;

wire n76,n77,n78,n79,n80,n81,n82,n83,n84,
n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,
n95,n96,n97,n98,n99,n100,n101,n102,n103,n104,
n105,n106,n107,n108,n109,n110,n111,n112,n113,n114,
n115,n116,n117,n118,n119,n120,n121,n122,n123,n124,
n125,n126,n127,n128,n129,n130,n131,n132,n133,n134,
n135,n136,n137,n138,n139,n140,n141,n142,n143,n144,
n145,n146,n147,n148,n149,n150,n151,n152,n153,n154,
n155,n156,n157,n158,n159,n160,n161,n162,n163,n164,
n165,n166,n167,n168,n169,n170,n171,n172,n173,n174,
n175,n176,n177,n178,n179,n180,n181,n182,n183,n184,
n185,n186,n187,n188,n189,n190,n191,n192,n193,n194,
n195,n196,n197,n198,n199,n200,n201,n202,n203,n204,
n205,n206,n207,n208,n209,n210,n211,n212,n213,n214,
n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,
n225,n226,n227,n228,n229,n230,n231,n232,n233,n234,
n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,
n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,
n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,
n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,
n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,
n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,
n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,
n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,
n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,
n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,
n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,
n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,
n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,
n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,
n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,
n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,
n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,
n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,
n415,n416,n417,n418,n419,n420,n421,n422,n423,n424,
n425,n426,n427,n428,n429,n431,n432,n433,n434,n435,
n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,
n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,
n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,
n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,
n476,n477,n478,n479,n480,n481,n482,n483,n484,n485,
n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,
n496,n497,n498,n499,n500,n501,n502,n503,n504,n505,
n506,n507,n508,n509,n510,n511,n512,n513,n514,n515,
n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,
n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,
n536,n537,n538,n539,n540,n541,n542,n543,n544,n545,
n546,n547,n548,n549,n550,n551,n552,n553,n554,n555,
n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,
n566,n567,n568,n569,n570,n571,n572,n573,n574,n575,
n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,
n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,
n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,
n606,n607,n608,n609,n610,n611,n612,n614,n615,n616,
n617,n618,n619,n620,n621,n622,n623,n624,n625,n626,
n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,
n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,
n647,n648,n649,n650,n651,n652,n653,n654,n655,n656,
n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,
n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,
n677,n678,n679,n680,n681,n682,n683,n684,n685,n686,
n687,n688,n689,n690,n691,n692,n693,n694,n695,n696,
n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,
n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,
n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,
n727,n728,n729,n730,n731,n732,n733,n734,n735,n736,
n737,n738,n739,n740,n741,n742,n743,n744,n745,n746,
n747,n748,n749,n750,n751,n752,n753,n754,n755,n757,
n758,n759,n760,n761,n762,n763,n764,n765,n766,n767,
n768,n769,n770,n771,n772,n773,n774,n775,n776,n777,
n778,n779,n780,n781,n782,n783,n784,n785,n786,n787,
n788,n789,n790,n791,n792,n793,n794,n795,n796,n797,
n798,n799,n800,n801,n802,n803,n804,n805,n806,n807,
n808,n809,n810,n811,n812,n813,n814,n815,n816,n817,
n818,n819,n820,n821,n822,n823,n824,n825,n826,n827,
n828,n829,n830,n831,n832,n833,n834,n835,n836,n837,
n838,n839,n840,n841,n842,n843,n844,n845,n846,n847,
n848,n849,n850,n851,n852,n853,n854,n855,n856,n857,
n858,n859,n860,n861,n862,n863,n864,n865,n866,n867,
n868,n869,n870,n871,n872,n873,n874,n875,n876,n877,
n878,n879,n880,n881,n882,n883,n884,n885,n886,n887,
n888,n889,n890,n891,n892,n893,n894,n895,n896,n897,
n898,n899,n900,n901,n902,n903,n904,n905,n906,n907,
n908,n909,n910,n911,n912,n913,n914,n915,n916,n917,
n918,n919,n920,n921,n922,n923,n924,n925,n926,n927,
n928,n929,n930,n931,n932,n933,n934,n935,n936,n937,
n938,n939,n940,n941,n942,n943,n944,n945,n946,n947,
n948,n949,n950,n951,n952,n953,n954,n955,n956,n957,
n958,n959,n960,n961,n962,n963,n964,n965,n966,n967,
n968,n969,n970,n971,n972,n973,n974,n975,n976,n977,
n978,n979,n980,n981,n982,n983,n984,n985,n986,n987,
n988,n989,n990,n991,n992,n993,n994,n995,n996,n997,
n998,n999,n1000,n1001,n1002,n1003,n1004,n1005,n1006,n1007,
n1008,n1009,n1010,n1011,n1012,n1013,n1014,n1015,n1016,n1017,
n1018,n1019,n1020,n1021,n1022,n1023,n1024,n1025,n1026,n1027,
n1028,n1029,n1030,n1031,n1032,n1033,n1034,n1035,n1036,n1037,
n1038,n1039,n1040,n1041,n1042,n1043,n1044,n1045,n1046,n1047,
n1048,n1049,n1050,n1051,n1052,n1053,n1054,n1055,n1056,n1057,
n1058,n1059,n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,
n1069,n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,
n1079,n1080,n1081,n1082,n1083,n1084,n1085,n1086,n1087,n1088,
n1089,n1090,n1091,n1092,n1093,n1094,n1095,n1096,n1097,n1098,
n1099,n1100,n1101,n1102,n1103,n1104,n1105,n1106,n1107,n1108,
n1109,n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,n1118,
n1119,n1120,n1121,n1122,n1123,n1124,n1125,n1126,n1127,n1128,
n1129,n1130,n1131,n1132,n1133,n1134,n1135,n1136,n1137,n1138,
n1139,n1140,n1141,n1142,n1143,n1144,n1145,n1146,n1147,n1148,
n1149,n1150,n1151,n1152,n1153,n1154,n1155,n1156,n1157,n1158,
n1159,n1160,n1161,n1162,n1163,n1164,n1165,n1166,n1167,n1168,
n1169,n1170,n1171,n1172,n1173,n1174,n1175,n1176,n1177,n1178,
n1179,n1180,n1181,n1182,n1183,n1184,n1185,n1186,n1187,n1188,
n1189,n1190,n1191,n1192,n1193,n1194,n1195,n1196,n1197,n1198,
n1199,n1200,n1201,n1202,n1203,n1204,n1205,n1206,n1207,n1208,
n1209,n1210,n1211,n1212,n1213,n1214,n1215,n1216,n1217,n1218,
n1219,n1220,n1221,n1222,n1223,n1224,n1225,n1226,n1227,n1228,
n1229,n1230,n1231,n1232,n1233,n1234,n1235,n1237,n1238,n1239,
n1240,n1241,n1242,n1243,n1244,n1245,n1246,n1247,n1248,n1249,
n1250,n1251,n1252,n1253,n1254,n1255,n1256,n1257,n1258,n1259,
n1260,n1261,n1262,n1263,n1264,n1265,n1266,n1267,n1268,n1269,
n1270,n1271,n1272,n1273,n1274,n1275,n1276,n1277,n1278,n1279,
n1280,n1281,n1282,n1283,n1284,n1285,n1286,n1287,n1288,n1289,
n1290,n1291,n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,
n1300,n1301,n1302,n1303,n1304,n1305,n1306,n1307,n1308,n1309,
n1310,n1311,n1312,n1313,n1314,n1315,n1316,n1317,n1318,n1319,
n1320,n1321,n1322,n1323,n1324,n1325,n1326,n1327,n1328,n1329,
n1330,n1331,n1332,n1333,n1334,n1335,n1336,n1337,n1338,n1339,
n1340,n1341,n1342,n1343,n1344,n1345,n1346,n1347,n1348,n1349,
n1350,n1351,n1352,n1353,n1354,n1355,n1356,n1357,n1358,n1359,
n1360,n1361,n1362,n1363,n1364,n1365,n1366,n1367,n1368,n1369,
n1370,n1371,n1372,n1373,n1374,n1375,n1376,n1377,n1378,n1379,
n1380,n1381,n1382,n1383,n1384,n1385,n1386,n1387,n1388,n1389,
n1390,n1391,n1392,n1393,n1394,n1395,n1396,n1397,n1398,n1399,
n1400,n1401,n1402,n1403,n1404,n1405,n1406,n1407,n1408,n1409,
n1410,n1411,n1412,n1413,n1414,n1415,n1416,n1417,n1418,n1419,
n1420,n1421,n1422,n1423,n1424,n1425,n1426,n1427,n1428,n1429,
n1430,n1431,n1432,n1433,n1434,n1435,n1436,n1437,n1438,n1439,
n1440,n1441,n1442,n1443,n1444,n1445,n1446,n1447,n1448,n1449,
n1450,n1451,n1452,n1453,n1454,n1455,n1456,n1457,n1458,n1459,
n1460,n1461,n1462,n1463,n1464,n1465,n1466,n1467,n1468,n1469,
n1470,n1471,n1472,n1473,n1474,n1475,n1476,n1477,n1478,n1479,
n1480,n1481,n1482,n1483,n1484,n1485,n1486,n1487,n1488,n1489,
n1490,n1491,n1492,n1493,n1494,n1495,n1496,n1497,n1498,n1499,
n1500,n1501,n1502,n1503,n1504,n1505,n1506,n1507,n1509,n1510,
n1511,n1512,n1513,n1514,n1515,n1516,n1517,n1518,n1519,n1520,
n1521,n1522,n1523,n1524,n1525,n1526,n1527,n1528,n1529,n1530,
n1531,n1532,n1533,n1534,n1535,n1536,n1537,n1538,n1539,n1540,
n1541,n1542,n1543,n1544,n1545,n1546,n1547,n1548,n1549,n1550,
n1551,n1552,n1553,n1554,n1555,n1556,n1557,n1558,n1559,n1560,
n1561,n1562,n1563,n1564,n1565,n1566,n1567,n1568,n1569,n1570,
n1571,n1572,n1573,n1574,n1575,n1576,n1577,n1578,n1579,n1580,
n1581,n1582,n1583,n1584,n1585,n1586,n1587,n1588,n1589,n1590,
n1591,n1592,n1593,n1594,n1595,n1596,n1597,n1598,n1599,n1600,
n1601,n1602,n1603,n1604,n1605,n1606,n1607,n1608,n1609,n1610,
n1611,n1612,n1613,n1614,n1615,n1616,n1617,n1618,n1619,n1620,
n1621,n1622,n1623,n1624,n1625,n1626,n1627,n1628,n1629,n1630,
n1631,n1632,n1633,n1634,n1635,n1636,n1637,n1638,n1639,n1640,
n1641,n1642,n1643,n1644,n1645,n1646,n1647,n1648,n1649,n1650,
n1651,n1652,n1653,n1654,n1655,n1656,n1657,n1658,n1659,n1660,
n1661,n1662,n1663,n1664,n1665,n1666,n1667,n1668,n1669,n1670,
n1671,n1672,n1673,n1674,n1675,n1676,n1677,n1678,n1679,n1680,
n1681,n1682,n1683,n1684,n1685,n1686,n1687,n1688,n1689,n1690,
n1692,n1693,n1694,n1695,n1696,n1697,n1698,n1699,n1700,n1701,
n1702,n1703,n1704,n1705,n1706,n1707,n1708,n1709,n1710,n1711,
n1712,n1713,n1714,n1715,n1716,n1717,n1718,n1719,n1720,n1721,
n1722,n1723,n1724,n1725,n1726,n1727,n1728,n1729,n1730,n1731,
n1732,n1733,n1734,n1735,n1736,n1737,n1738,n1739,n1740,n1741,
n1742,n1743,n1744,n1745,n1746,n1747,n1748,n1749,n1750,n1751,
n1752,n1753,n1754,n1755,n1756,n1757,n1758,n1759,n1760,n1761,
n1762,n1763,n1764,n1765,n1766,n1767,n1768,n1769,n1770,n1771,
n1772,n1773,n1774,n1775,n1776,n1777,n1778,n1779,n1780,n1781,
n1783,n1784,n1785,n1786,n1787,n1788,n1789,n1790,n1791,n1792,
n1793,n1794,n1795,n1796,n1797,n1798,n1800,n1801,n1802,n1803,
n1804,n1805,n1806,n1807,n1808,n1809,n1810,n1811,n1812,n1813,
n1814,n1815,n1816,n1817,n1818,n1819,n1820,n1821,n1822,n1823,
n1825,n1826,n1827,n1828,n1829,n1830,n1831,n1832,n1833,n1834,
n1835,n1836,n1837,n1838,n1839,n1840,n1841,n1842,n1843,n1844,
n1845,n1846,n1847,n1848,n1849,n1850,n1851,n1852,n1853,n1854,
n1856,n1857,n1858,n1859,n1860,n1861,n1862,n1863,n1864,n1865,
n1866,n1867,n1868,n1869,n1870,n1871,n1872,n1873,n1874,n1875,
n1876,n1877,n1878,n1879,n1880,n1881,n1882,n1883,n1885,n1886,
n1887,n1888,n1889,n1890,n1891,n1892,n1893,n1894,n1895,n1896,
n1897,n1898,n1899,n1900,n1901,n1902,n1904,n1905,n1906,n1907,
n1908,n1909,n1910,n1911,n1912,n1913,n1914,n1915,n1916,n1917,
n1919,n1920,n1921,n1922,n1923,n1924,n1925,n1926,n1927,n1928,
n1931,n1932,n1933,n1934,n1935,n1936,n1937,n1938,n1939,n1940,
n1941,n1942,n1943,n1944,n1945,n1946,n1947,n1948,n1949,n1950,
n1951,n1952,n1953,n1954,n1955,n1956,n1957,n1958,n1959,n1960,
n1961,n1962,n1963,n1964,n1965,n1966,n1967,n1968,n1969,n1970,
n1971,n1972,n1974,n1975,n1976,n1977,n1978,n1979,n1980,n1981,
n1982,n1983,n1984,n1985,n1986,n1987,n1988,n1989,n1990,n1991,
n1992,n1993,n1994,n1995,n1996,n1997,n1998,n1999,n2000,n2001,
n2002,n2003,n2004,n2005,n2006,n2007,n2008,n2009,n2010,n2011,
n2012,n2013,n2014,n2015,n2016,n2017,n2018,n2019,n2020,n2021,
n2022,n2023,n2024,n2025,n2026,n2027,n2028,n2029,n2030,n2031,
n2032,n2033,n2034,n2035,n2036,n2037,n2038,n2039,n2040,n2041,
n2042,n2043,n2044,n2045,n2046,n2047,n2048,n2049,n2050,n2051,
n2052,n2053,n2054,n2055,n2056,n2057,n2058,n2059,n2060,n2061,
n2062,n2063,n2064,n2065,n2066,n2067,n2068,n2069,n2070,n2071,
n2072,n2073,n2074,n2075,n2076,n2077,n2078,n2079,n2080,n2081,
n2082,n2083,n2084,n2085,n2086,n2087,n2088,n2089,n2090,n2091,
n2092,n2093,n2094,n2095,n2096,n2097,n2098,n2099,n2100,n2101,
n2102,n2103,n2104,n2105,n2106,n2107,n2108,n2109,n2110,n2111,
n2112,n2113,n2114,n2115,n2116,n2117,n2118,n2119,n2120,n2121,
n2122,n2123,n2124,n2125,n2126,n2128,n2129,n2130,n2131,n2132,
n2133,n2134,n2135,n2136,n2137,n2138,n2139,n2140,n2141,n2142,
n2143,n2144,n2145,n2146,n2147,n2148,n2149,n2150,n2151,n2152,
n2153,n2154,n2155,n2156,n2157,n2158,n2159,n2160,n2161,n2162,
n2163,n2164,n2165,n2166,n2167,n2168,n2169,n2170,n2171,n2172,
n2173,n2174,n2175,n2176,n2177,n2178,n2179,n2180,n2181,n2182,
n2183,n2184,n2185,n2186,n2187,n2188,n2189,n2190,n2191,n2192,
n2193,n2194,n2195,n2196,n2197,n2198,n2199,n2200,n2201,n2202,
n2203,n2204,n2205,n2206,n2207,n2208,n2209,n2210,n2211,n2212,
n2213,n2214,n2215,n2216,n2217,n2218,n2219,n2220,n2221,n2222,
n2223,n2224,n2225,n2226,n2227,n2228,n2229,n2230,n2231,n2232,
n2233,n2234,n2235,n2236,n2237,n2238,n2239,n2240,n2241,n2242,
n2243,n2244,n2245,n2246,n2247,n2248,n2249,n2250,n2251,n2252,
n2253,n2254,n2255,n2256,n2257,n2258,n2259,n2260,n2261,n2262,
n2263,n2264,n2265,n2266,n2267,n2268,n2269,n2270,n2271,n2272,
n2273,n2274,n2275,n2276,n2277,n2278,n2279,n2280,n2281,n2282,
n2283,n2284,n2285,n2286,n2287,n2288,n2289,n2290,n2291,n2292,
n2293,n2294,n2295,n2296,n2297,n2298,n2299,n2301,n2302,n2303,
n2304,n2305,n2306,n2307,n2308,n2309,n2310,n2311,n2312,n2313,
n2314,n2315,n2316,n2317,n2318,n2319,n2320,n2321,n2322,n2323,
n2324,n2325,n2326,n2327,n2328,n2329,n2330,n2331,n2332,n2333,
n2334,n2335,n2336,n2337,n2338,n2339,n2340,n2341,n2342,n2343,
n2344,n2345,n2346,n2347,n2348,n2349,n2350,n2351,n2352,n2353,
n2354,n2355,n2356,n2357,n2358,n2359,n2361,n2362,n2363,n2364,
n2365,n2366,n2367,n2368,n2369,n2370,n2371,n2372,n2373,n2374,
n2375,n2376,n2377,n2378,n2379,n2380,n2381,n2382,n2383,n2384,
n2385,n2386,n2387,n2388,n2389,n2390,n2391,n2392,n2393,n2394,
n2395,n2396,n2397,n2398,n2399,n2400,n2401,n2402,n2403,n2404,
n2405,n2406,n2407,n2408,n2409,n2410,n2411,n2412,n2413,n2414,
n2415,n2416,n2417,n2418,n2419,n2420,n2421,n2422,n2423,n2424,
n2425,n2426,n2427,n2428,n2429,n2430,n2431,n2432,n2433,n2434,
n2435,n2436,n2437,n2438,n2439,n2440,n2441,n2442,n2443,n2444,
n2445,n2446,n2447,n2448,n2449,n2450,n2451,n2452,n2453,n2454,
n2455,n2456,n2457,n2458,n2459,n2460,n2461,n2462,n2463,n2464,
n2465,n2466,n2467,n2468,n2469,n2470,n2471,n2472,n2473,n2474,
n2475,n2476,n2477,n2478,n2479,n2480,n2481,n2482,n2483,n2484,
n2485,n2486,n2487,n2488,n2489,n2490,n2492,n2493,n2494,n2495,
n2496,n2497,n2498,n2499,n2500,n2501,n2502,n2503,n2504,n2505,
n2506,n2507,n2508,n2509,n2510,n2511,n2512,n2513,n2514,n2515,
n2516,n2517,n2518,n2519,n2520,n2521,n2522,n2523,n2524,n2525,
n2526,n2527,n2528,n2529,n2530,n2531,n2532,n2533,n2534,n2535,
n2536,n2537,n2538,n2539,n2540,n2541,n2542,n2543,n2544,n2545,
n2546,n2547,n2548,n2549,n2550,n2551,n2552,n2554,n2555,n2556,
n2557,n2558,n2559,n2560,n2561,n2562,n2563,n2564,n2565,n2566,
n2567,n2568,n2569,n2570,n2571,n2572,n2573,n2574,n2575,n2576,
n2577,n2578,n2579,n2580,n2581,n2582,n2583,n2584,n2585,n2586,
n2587,n2588,n2589,n2590,n2591,n2592,n2593,n2594,n2595,n2596,
n2597,n2598,n2599,n2600,n2601,n2602,n2603,n2604,n2605,n2606,
n2607,n2608,n2609,n2610,n2611,n2612,n2613,n2614,n2615,n2616,
n2618,n2619,n2620,n2621,n2622,n2623,n2624,n2625,n2626,n2627,
n2628,n2629,n2630,n2631,n2632,n2633,n2634,n2635,n2636,n2637,
n2638,n2639,n2640,n2641,n2642,n2643,n2644,n2645,n2646,n2647,
n2648,n2649,n2650,n2651,n2652,n2653,n2654,n2655,n2656,n2657,
n2658,n2659,n2660,n2661,n2662,n2663,n2664,n2665,n2666,n2667,
n2668,n2669,n2670,n2671,n2672,n2673,n2674,n2675,n2676,n2677,
n2678,n2679,n2680,n2681,n2682,n2683,n2684,n2685,n2686,n2687,
n2688,n2689,n2690,n2691,n2692,n2693,n2694,n2695,n2696,n2697,
n2698,n2699,n2700,n2701,n2702,n2703,n2704,n2705,n2706,n2707,
n2708,n2709,n2710,n2711,n2712,n2713,n2714,n2715,n2716,n2717,
n2718,n2719,n2720,n2721,n2722,n2723,n2724,n2725,n2726,n2727,
n2728,n2729,n2730,n2731,n2732,n2733,n2734,n2735,n2736,n2737,
n2738,n2739,n2740,n2741,n2742,n2743,n2744,n2745,n2746,n2747,
n2748,n2749,n2750,n2751,n2752,n2753,n2754,n2755,n2756,n2757,
n2758,n2759,n2760,n2761,n2762,n2763,n2764,n2765,n2766,n2767,
n2768,n2769,n2771,n2772,n2773,n2774,n2775,n2776,n2777,n2778,
n2779,n2780,n2781,n2782,n2783,n2784,n2785,n2786,n2787,n2788,
n2789,n2790,n2791,n2792,n2793,n2794,n2795,n2796,n2797,n2798,
n2799,n2800,n2801,n2802,n2803,n2804,n2805,n2806,n2807,n2808,
n2809,n2810,n2811,n2812,n2813,n2814,n2815,n2816,n2817,n2818,
n2819,n2820,n2821,n2822,n2823,n2824,n2825,n2826,n2827,n2828,
n2829,n2830,n2831,n2832,n2833,n2834,n2835,n2836,n2837,n2838,
n2839,n2840,n2841,n2842,n2843,n2844,n2845,n2846,n2847,n2848,
n2849,n2850,n2851,n2852,n2853,n2854,n2855,n2856,n2857,n2858,
n2859,n2860,n2861,n2862,n2863,n2864,n2865,n2866,n2867,n2868,
n2869,n2870,n2871,n2872,n2873,n2874,n2875,n2876,n2877,n2878,
n2879,n2880,n2881,n2882,n2883,n2884,n2885,n2886,n2887,n2888,
n2889,n2890,n2891,n2892,n2894,n2895,n2896,n2897,n2898,n2899,
n2900,n2901,n2902,n2903,n2904,n2905,n2906,n2907,n2908,n2909,
n2910,n2911,n2912,n2913,n2914,n2915,n2916,n2917,n2918,n2919,
n2920,n2921,n2922,n2923,n2924,n2925,n2926,n2927,n2928,n2929,
n2930,n2931,n2932,n2933,n2934,n2935,n2936,n2937,n2938,n2939,
n2940,n2941,n2942,n2943,n2944,n2945,n2946,n2947,n2948,n2949,
n2950,n2951,n2952,n2953,n2954,n2955,n2956,n2957,n2958,n2959,
n2960,n2961,n2962,n2963,n2964,n2965,n2966,n2967,n2968,n2969,
n2970,n2971,n2972,n2973,n2974,n2975,n2976,n2977,n2978,n2979,
n2980,n2981,n2982,n2983,n2984,n2985,n2986,n2987,n2988,n2989,
n2990,n2991,n2992,n2993,n2994,n2995,n2996,n2997,n2998,n2999,
n3000,n3001,n3003,n3004,n3005,n3006,n3007,n3008,n3009,n3010,
n3011,n3012,n3013,n3014,n3015,n3016,n3017,n3018,n3019,n3020,
n3021,n3022,n3023,n3024,n3025,n3026,n3027,n3028,n3030,n3031,
n3032,n3033,n3034,n3035,n3036,n3037,n3038,n3039,n3040,n3041,
n3042,n3043,n3044,n3045,n3046,n3047,n3048,n3049,n3050,n3051,
n3052,n3053,n3054,n3055,n3056,n3057,n3058,n3059,n3060,n3061,
n3062,n3063,n3064,n3065,n3066,n3067,n3068,n3069,n3070,n3071,
n3072,n3073,n3074,n3075,n3076,n3077,n3078,n3079,n3080,n3081,
n3082,n3083,n3084,n3085,n3087,n3088,n3089,n3090,n3091,n3092,
n3093,n3094,n3095,n3096,n3097,n3098,n3099,n3101,n3102,n3103,
n3104,n3105,n3106,n3107,n3108,n3109,n3110,n3111,n3112,n3113,
n3114,n3115,n3116,n3117,n3118,n3119,n3120,n3121,n3122,n3123,
n3124,n3125,n3126,n3127,n3128,n3129,n3130,n3131,n3132,n3133,
n3134,n3136,n3137,n3138,n3139,n3140,n3141,n3142,n3143,n3144,
n3145,n3146,n3147,n3148,n3149,n3150,n3151,n3152,n3153,n3154,
n3155,n3156,n3157,n3158,n3159,n3160,n3161,n3162,n3163,n3164,
n3165,n3166,n3167,n3168,n3169,n3170,n3172,n3173,n3174,n3175,
n3176,n3177,n3178,n3179,n3180,n3181,n3182,n3183,n3184,n3185,
n3186,n3187,n3188,n3189,n3190,n3191,n3192,n3193,n3194,n3195,
n3196,n3197,n3198,n3199,n3200,n3201,n3202,n3203,n3204,n3205,
n3206,n3207,n3208,n3209,n3210,n3211,n3213,n3214,n3216,n3217,
n3218,n3219,n3220,n3221,n3222,n3223,n3224,n3225,n3226,n3227,
n3228,n3229,n3230,n3231,n3232,n3233,n3234,n3235,n3236,n3237,
n3238,n3239,n3240,n3241,n3242,n3243,n3244,n3245,n3246,n3247,
n3248,n3249,n3250,n3251,n3252,n3253,n3254,n3255,n3256,n3257,
n3258,n3259,n3260,n3261,n3262,n3263,n3264,n3265,n3266,n3267,
n3268,n3269,n3270,n3271,n3272,n3273,n3274,n3275,n3276,n3277,
n3278,n3279,n3280,n3281,n3282,n3283,n3284,n3285,n3286,n3287,
n3288,n3289,n3290,n3291,n3292,n3293,n3294,n3295,n3296,n3297,
n3298,n3299,n3300,n3301,n3302,n3303,n3304,n3305,n3306,n3307,
n3308,n3309,n3310,n3311,n3312,n3313,n3314,n3315,n3316,n3317,
n3318,n3319,n3320,n3321,n3322,n3323,n3324,n3325,n3326,n3327,
n3328,n3329,n3330,n3331,n3332,n3333,n3334,n3335,n3336,n3337,
n3338,n3339,n3340,n3341,n3342,n3343,n3344,n3345,n3346,n3347,
n3348,n3349,n3350,n3351,n3352,n3353,n3354,n3355,n3356,n3357,
n3358,n3359,n3360,n3361,n3362,n3363,n3364,n3365,n3366,n3367,
n3368,n3369,n3370,n3371,n3372,n3373,n3374,n3375,n3376,n3377,
n3378,n3379,n3380,n3381,n3382,n3383,n3384,n3385,n3386,n3387,
n3388,n3389,n3390,n3391,n3392,n3393,n3394,n3395,n3396,n3397,
n3398,n3399,n3400,n3401,n3402,n3403,n3404,n3405,n3406,n3407,
n3408,n3409,n3410,n3411,n3412,n3413,n3414,n3415,n3416,n3417,
n3419,n3420,n3421,n3422,n3423,n3424,n3425,n3426,n3427,n3428,
n3429,n3430,n3431,n3432,n3433,n3434,n3435,n3436,n3437,n3438,
n3439,n3440,n3441,n3442,n3443,n3444,n3445,n3446,n3447,n3448,
n3449,n3450,n3451,n3452,n3453,n3454,n3455,n3456,n3457,n3458,
n3459,n3460,n3461,n3462,n3463,n3464,n3465,n3466,n3467,n3468,
n3469,n3470,n3471,n3472,n3473,n3474,n3475,n3476,n3477,n3478,
n3479,n3480,n3481,n3482,n3483,n3484,n3485,n3486,n3487,n3488,
n3489,n3490,n3491,n3492,n3493,n3494,n3495,n3496,n3497,n3498,
n3499,n3500,n3501,n3502,n3503,n3504,n3505,n3506,n3507,n3508,
n3509,n3510,n3511,n3512,n3513,n3514,n3515,n3516,n3517,n3518,
n3519,n3520,n3521,n3522,n3523,n3524,n3525,n3526,n3527,n3528,
n3529,n3530,n3531,n3532,n3533,n3534,n3535,n3536,n3537,n3538,
n3539,n3540,n3541,n3542,n3543,n3544,n3545,n3546,n3547,n3548,
n3549,n3550,n3551,n3552,n3553,n3554,n3555,n3556,n3557,n3558,
n3559,n3560,n3561,n3562,n3563,n3564,n3565,n3566,n3567,n3568,
n3569,n3570,n3571,n3572,n3573,n3574,n3575,n3576,n3577,n3578,
n3579,n3580,n3581,n3582,n3583,n3584,n3585,n3586,n3587,n3588,
n3589,n3590,n3591,n3592,n3593;
not gate_0(n76,pi00);
not gate_1(n77,pi01);
not gate_2(n78,pi02);
not gate_3(n79,pi03);
not gate_4(n80,pi04);
not gate_5(n81,pi05);
not gate_6(n82,pi06);
not gate_7(n83,pi07);
not gate_8(n84,pi09);
not gate_9(n85,pi11);
not gate_10(n86,pi12);
not gate_11(n87,pi13);
not gate_12(n88,pi14);
not gate_13(n89,pi15);
not gate_14(n90,pi16);
not gate_15(n91,pi17);
not gate_16(n92,pi18);
not gate_17(n93,pi19);
not gate_18(n94,pi20);
not gate_19(n95,pi21);
not gate_20(n96,pi22);
not gate_21(n97,pi23);
not gate_22(n98,pi24);
not gate_23(n99,pi25);
not gate_24(n100,pi26);
not gate_25(n101,pi28);
not gate_26(n102,pi29);
not gate_27(n103,pi30);
not gate_28(n104,pi31);
not gate_29(n105,pi32);
not gate_30(n106,pi33);
not gate_31(n107,pi34);
not gate_32(n108,pi35);
not gate_33(n109,pi36);
not gate_34(n110,pi37);
not gate_35(n111,pi38);
not gate_36(n112,pi39);
not gate_37(n113,pi40);
and gate_38(n114,pi02,n79);
not gate_39(n115,n114);
and gate_40(n116,pi04,n115);
not gate_41(n117,n116);
and gate_42(n118,pi35,pi37);
not gate_43(n119,n118);
and gate_44(n120,n117,n118);
and gate_45(n121,n77,n120);
not gate_46(n122,n121);
and gate_47(n123,n77,n78);
and gate_48(n124,n79,n80);
and gate_49(n125,n123,n124);
not gate_50(n126,n125);
and gate_51(n127,n108,n126);
and gate_52(n128,n110,pi39);
not gate_53(n129,n128);
and gate_54(n130,pi37,n112);
not gate_55(n131,n130);
and gate_56(n132,n129,n131);
not gate_57(n133,n132);
and gate_58(n134,pi40,n133);
not gate_59(n135,n134);
and gate_60(n136,n127,n134);
not gate_61(n137,n136);
and gate_62(n138,n122,n137);
not gate_63(n139,n138);
and gate_64(n140,pi38,n139);
not gate_65(n141,n140);
and gate_66(n142,pi01,n78);
and gate_67(n143,n79,pi04);
and gate_68(n144,n142,n143);
not gate_69(n145,n144);
and gate_70(n146,n111,n145);
and gate_71(n147,pi37,n113);
not gate_72(n148,n147);
and gate_73(n149,n146,n147);
and gate_74(n150,pi35,n149);
not gate_75(n151,n150);
and gate_76(n152,n141,n151);
not gate_77(n153,n152);
and gate_78(n154,pi36,n153);
not gate_79(n155,n154);
and gate_80(n156,n109,pi37);
not gate_81(n157,n156);
and gate_82(n158,pi35,n156);
and gate_83(n159,pi39,n113);
not gate_84(n160,n159);
and gate_85(n161,pi38,n159);
and gate_86(n162,n158,n161);
not gate_87(n163,n162);
and gate_88(n164,n155,n163);
not gate_89(n165,n164);
and gate_90(n166,n107,n165);
not gate_91(n167,n166);
and gate_92(n168,n110,n111);
not gate_93(n169,n168);
and gate_94(n170,n108,n109);
and gate_95(n171,n168,n170);
not gate_96(n172,n171);
and gate_97(n173,n117,n171);
and gate_98(n174,pi34,n173);
and gate_99(n175,n77,n174);
not gate_100(n176,n175);
and gate_101(n177,n167,n176);
not gate_102(n178,n177);
and gate_103(n179,pi00,n178);
not gate_104(n180,n179);
and gate_105(n181,pi38,pi39);
not gate_106(n182,n181);
and gate_107(n183,n110,n181);
not gate_108(n184,n183);
and gate_109(n185,n111,n112);
not gate_110(n186,n185);
and gate_111(n187,pi37,n185);
not gate_112(n188,n187);
and gate_113(n189,n184,n188);
not gate_114(n190,n189);
and gate_115(n191,n126,n190);
not gate_116(n192,n191);
and gate_117(n193,pi38,n112);
not gate_118(n194,n193);
and gate_119(n195,n85,n86);
not gate_120(n196,n195);
and gate_121(n197,pi15,n196);
not gate_122(n198,n197);
and gate_123(n199,n87,n198);
not gate_124(n200,n199);
and gate_125(n201,n81,n200);
not gate_126(n202,n201);
and gate_127(n203,pi37,n202);
not gate_128(n204,n203);
and gate_129(n205,n111,pi39);
not gate_130(n206,n205);
and gate_131(n207,n204,n205);
not gate_132(n208,n207);
and gate_133(n209,n194,n208);
not gate_134(n210,n209);
and gate_135(n211,pi40,n210);
not gate_136(n212,n211);
and gate_137(n213,n192,n212);
not gate_138(n214,n213);
and gate_139(n215,pi34,n214);
not gate_140(n216,n215);
and gate_141(n217,n112,pi40);
not gate_142(n218,n217);
and gate_143(n219,pi38,n217);
not gate_144(n220,n219);
and gate_145(n221,n107,pi37);
and gate_146(n222,n111,n159);
not gate_147(n223,n222);
and gate_148(n224,n221,n222);
not gate_149(n225,n224);
and gate_150(n226,n220,n225);
not gate_151(n227,n226);
and gate_152(n228,pi29,pi30);
and gate_153(n229,n101,n228);
not gate_154(n230,n229);
and gate_155(n231,n102,n103);
not gate_156(n232,n231);
and gate_157(n233,pi28,n231);
not gate_158(n234,n233);
and gate_159(n235,n230,n234);
not gate_160(n236,n235);
and gate_161(n237,n227,n236);
not gate_162(n238,n237);
and gate_163(n239,n86,pi13);
not gate_164(n240,n239);
and gate_165(n241,n112,n240);
not gate_166(n242,n241);
and gate_167(n243,n85,n242);
not gate_168(n244,n243);
and gate_169(n245,pi12,pi15);
not gate_170(n246,n245);
and gate_171(n247,pi13,n89);
not gate_172(n248,n247);
and gate_173(n249,n112,n248);
not gate_174(n250,n249);
and gate_175(n251,n246,n250);
not gate_176(n252,n251);
and gate_177(n253,n244,n252);
and gate_178(n254,n84,n90);
not gate_179(n255,n254);
and gate_180(n256,n197,n254);
not gate_181(n257,n256);
and gate_182(n258,n253,n257);
not gate_183(n259,n258);
and gate_184(n260,n113,n259);
not gate_185(n261,n260);
and gate_186(n262,n90,n91);
not gate_187(n263,n262);
and gate_188(n264,pi39,n196);
and gate_189(n265,pi12,n113);
not gate_190(n266,n265);
and gate_191(n267,n264,n266);
and gate_192(n268,n262,n267);
and gate_193(n269,pi15,n268);
not gate_194(n270,n269);
and gate_195(n271,n261,n270);
not gate_196(n272,n271);
and gate_197(n273,n110,n272);
not gate_198(n274,n273);
and gate_199(n275,n110,pi40);
not gate_200(n276,n275);
and gate_201(n277,pi16,pi17);
not gate_202(n278,n277);
and gate_203(n279,n197,n278);
not gate_204(n280,n279);
and gate_205(n281,n275,n280);
not gate_206(n282,n281);
and gate_207(n283,pi39,n282);
and gate_208(n284,n84,n283);
not gate_209(n285,n284);
and gate_210(n286,n274,n285);
not gate_211(n287,n286);
and gate_212(n288,pi38,n287);
not gate_213(n289,n288);
and gate_214(n290,n113,n131);
not gate_215(n291,n290);
and gate_216(n292,n111,n291);
not gate_217(n293,n292);
and gate_218(n294,n129,n293);
not gate_219(n295,n294);
and gate_220(n296,pi13,n198);
not gate_221(n297,n296);
and gate_222(n298,n257,n297);
not gate_223(n299,n298);
and gate_224(n300,n295,n299);
not gate_225(n301,n300);
and gate_226(n302,pi09,pi16);
not gate_227(n303,n302);
and gate_228(n304,n196,n303);
and gate_229(n305,n187,n304);
and gate_230(n306,n91,n305);
and gate_231(n307,pi15,n306);
not gate_232(n308,n307);
and gate_233(n309,n301,n308);
and gate_234(n310,n289,n309);
not gate_235(n311,n310);
and gate_236(n312,n107,n311);
not gate_237(n313,n312);
and gate_238(n314,n238,n313);
not gate_239(n315,n314);
and gate_240(n316,n104,n315);
and gate_241(n317,n81,n316);
not gate_242(n318,n317);
and gate_243(n319,n216,n318);
not gate_244(n320,n319);
and gate_245(n321,n108,n320);
not gate_246(n322,n321);
and gate_247(n323,n182,n186);
not gate_248(n324,n323);
and gate_249(n325,n198,n324);
not gate_250(n326,n325);
and gate_251(n327,n112,n113);
not gate_252(n328,n327);
and gate_253(n329,n111,n327);
not gate_254(n330,n329);
and gate_255(n331,n326,n330);
not gate_256(n332,n331);
and gate_257(n333,pi13,n332);
not gate_258(n334,n333);
and gate_259(n335,pi24,pi40);
not gate_260(n336,n335);
and gate_261(n337,n324,n336);
not gate_262(n338,n337);
and gate_263(n339,n84,n92);
not gate_264(n340,n339);
and gate_265(n341,n95,pi22);
and gate_266(n342,n340,n341);
not gate_267(n343,n342);
and gate_268(n344,n181,n343);
not gate_269(n345,n344);
and gate_270(n346,n338,n345);
not gate_271(n347,n346);
and gate_272(n348,n197,n347);
not gate_273(n349,n348);
and gate_274(n350,n334,n349);
not gate_275(n351,n350);
and gate_276(n352,n110,n351);
not gate_277(n353,n352);
and gate_278(n354,pi18,pi19);
not gate_279(n355,n354);
and gate_280(n356,n84,n355);
not gate_281(n357,n356);
and gate_282(n358,n92,n93);
not gate_283(n359,n358);
and gate_284(n360,pi23,n359);
and gate_285(n361,n357,n360);
not gate_286(n362,n361);
and gate_287(n363,n341,n361);
not gate_288(n364,n363);
and gate_289(n365,pi37,n364);
not gate_290(n366,n365);
and gate_291(n367,pi24,n366);
not gate_292(n368,n367);
and gate_293(n369,n197,n368);
not gate_294(n370,n369);
and gate_295(n371,n297,n370);
not gate_296(n372,n371);
and gate_297(n373,n111,n217);
not gate_298(n374,n373);
and gate_299(n375,n372,n373);
not gate_300(n376,n375);
and gate_301(n377,n353,n376);
not gate_302(n378,n377);
and gate_303(n379,n107,pi35);
and gate_304(n380,n378,n379);
and gate_305(n381,n81,n380);
not gate_306(n382,n381);
and gate_307(n383,n322,n382);
not gate_308(n384,n383);
and gate_309(n385,n109,n384);
not gate_310(n386,n385);
and gate_311(n387,n99,n100);
not gate_312(n388,n387);
and gate_313(n389,n110,n112);
not gate_314(n390,n389);
and gate_315(n391,n387,n389);
not gate_316(n392,n391);
and gate_317(n393,pi37,n159);
not gate_318(n394,n393);
and gate_319(n395,n392,n394);
not gate_320(n396,n395);
and gate_321(n397,pi35,n396);
not gate_322(n398,n397);
and gate_323(n399,pi11,n108);
and gate_324(n400,pi39,pi40);
not gate_325(n401,n400);
and gate_326(n402,n110,n400);
not gate_327(n403,n402);
and gate_328(n404,n399,n402);
not gate_329(n405,n404);
and gate_330(n406,n398,n405);
not gate_331(n407,n406);
and gate_332(n408,n111,n407);
not gate_333(n409,n408);
and gate_334(n410,pi38,n113);
not gate_335(n411,n410);
and gate_336(n412,pi10,pi27);
not gate_337(n413,n412);
and gate_338(n414,n112,n413);
not gate_339(n415,n414);
and gate_340(n416,n132,n415);
and gate_341(n417,n410,n416);
and gate_342(n418,n108,n417);
not gate_343(n419,n418);
and gate_344(n420,n409,n419);
not gate_345(n421,n420);
and gate_346(n422,n107,pi36);
and gate_347(n423,n421,n422);
not gate_348(n424,n423);
and gate_349(n425,n386,n424);
and gate_350(n426,n180,n425);
not gate_351(n427,n426);
and gate_352(n428,n83,n105);
and gate_353(n429,pi33,n428);
and gate_354(po00,n427,n429);
and gate_355(n431,n84,n278);
not gate_356(n432,n431);
and gate_357(n433,pi15,n263);
and gate_358(n434,pi12,n433);
and gate_359(n435,n187,n434);
and gate_360(n436,n432,n435);
not gate_361(n437,n436);
and gate_362(n438,pi31,n437);
not gate_363(n439,n438);
and gate_364(n440,pi09,n263);
not gate_365(n441,n440);
and gate_366(n442,n278,n441);
not gate_367(n443,n442);
and gate_368(n444,n86,pi37);
and gate_369(n445,n185,n444);
not gate_370(n446,n445);
and gate_371(n447,n110,pi38);
not gate_372(n448,n447);
and gate_373(n449,n400,n447);
not gate_374(n450,n449);
and gate_375(n451,n446,n450);
not gate_376(n452,n451);
and gate_377(n453,pi11,n452);
not gate_378(n454,n453);
and gate_379(n455,pi11,pi14);
not gate_380(n456,n455);
and gate_381(n457,n187,n456);
not gate_382(n458,n457);
and gate_383(n459,n450,n458);
not gate_384(n460,n459);
and gate_385(n461,pi12,n460);
not gate_386(n462,n461);
and gate_387(n463,n454,n462);
not gate_388(n464,n463);
and gate_389(n465,n443,n464);
and gate_390(n466,pi15,n465);
not gate_391(n467,n466);
and gate_392(n468,n111,n328);
not gate_393(n469,n468);
and gate_394(n470,n401,n469);
not gate_395(n471,n470);
and gate_396(n472,n110,n471);
not gate_397(n473,n472);
and gate_398(n474,n188,n473);
not gate_399(n475,n474);
and gate_400(n476,n199,n475);
not gate_401(n477,n476);
and gate_402(n478,n467,n477);
and gate_403(n479,n439,n478);
not gate_404(n480,n479);
and gate_405(n481,n108,n480);
not gate_406(n482,n481);
and gate_407(n483,n87,n325);
not gate_408(n484,n483);
and gate_409(n485,pi24,n196);
and gate_410(n486,pi15,n485);
not gate_411(n487,n486);
and gate_412(n488,n217,n486);
not gate_413(n489,n488);
and gate_414(n490,n484,n489);
not gate_415(n491,n490);
and gate_416(n492,n110,n491);
not gate_417(n493,n492);
and gate_418(n494,pi40,n198);
not gate_419(n495,n494);
and gate_420(n496,pi37,n111);
not gate_421(n497,n496);
and gate_422(n498,n494,n496);
and gate_423(n499,n87,n498);
not gate_424(n500,n499);
and gate_425(n501,n493,n500);
not gate_426(n502,n501);
and gate_427(n503,pi35,n502);
not gate_428(n504,n503);
and gate_429(n505,n482,n504);
not gate_430(n506,n505);
and gate_431(n507,n81,n506);
not gate_432(n508,n507);
and gate_433(n509,pi12,n108);
and gate_434(n510,pi14,pi15);
and gate_435(n511,n443,n447);
and gate_436(n512,n510,n511);
and gate_437(n513,n509,n512);
and gate_438(n514,pi11,n513);
not gate_439(n515,n514);
and gate_440(n516,n119,n515);
not gate_441(n517,n516);
and gate_442(n518,pi40,n517);
not gate_443(n519,n518);
and gate_444(n520,pi35,n496);
not gate_445(n521,n520);
and gate_446(n522,n519,n521);
not gate_447(n523,n522);
and gate_448(n524,pi39,n523);
not gate_449(n525,n524);
and gate_450(n526,pi38,n327);
not gate_451(n527,n526);
and gate_452(n528,n118,n526);
not gate_453(n529,n528);
and gate_454(n530,n525,n529);
and gate_455(n531,n508,n530);
not gate_456(n532,n531);
and gate_457(n533,n109,n532);
not gate_458(n534,n533);
and gate_459(n535,pi37,pi38);
and gate_460(n536,n108,n535);
not gate_461(n537,n536);
and gate_462(n538,n85,pi12);
not gate_463(n539,n538);
and gate_464(n540,n168,n538);
not gate_465(n541,n540);
and gate_466(n542,n537,n541);
not gate_467(n543,n542);
and gate_468(n544,pi39,n543);
and gate_469(n545,pi36,n544);
not gate_470(n546,n545);
and gate_471(n547,pi35,n110);
not gate_472(n548,n547);
and gate_473(n549,n193,n547);
not gate_474(n550,n549);
and gate_475(n551,n546,n550);
not gate_476(n552,n551);
and gate_477(n553,pi40,n552);
not gate_478(n554,n553);
and gate_479(n555,n112,n387);
not gate_480(n556,n555);
and gate_481(n557,pi36,n110);
and gate_482(n558,pi38,n160);
not gate_483(n559,n558);
and gate_484(n560,n557,n559);
not gate_485(n561,n560);
and gate_486(n562,n556,n560);
and gate_487(n563,pi35,n562);
not gate_488(n564,n563);
and gate_489(n565,n554,n564);
and gate_490(n566,n534,n565);
not gate_491(n567,n566);
and gate_492(n568,n107,n567);
not gate_493(n569,n568);
and gate_494(n570,n400,n496);
not gate_495(n571,n570);
and gate_496(n572,n327,n447);
not gate_497(n573,n572);
and gate_498(n574,n571,n573);
not gate_499(n575,n574);
and gate_500(n576,n199,n575);
not gate_501(n577,n576);
and gate_502(n578,pi31,n572);
not gate_503(n579,n578);
and gate_504(n580,n577,n579);
not gate_505(n581,n580);
and gate_506(n582,n81,n581);
not gate_507(n583,n582);
and gate_508(n584,n78,n79);
not gate_509(n585,n584);
and gate_510(n586,n77,n584);
and gate_511(n587,n80,n400);
and gate_512(n588,n586,n587);
not gate_513(n589,n588);
and gate_514(n590,n328,n589);
not gate_515(n591,n590);
and gate_516(n592,n447,n591);
and gate_517(n593,pi34,n592);
not gate_518(n594,n593);
and gate_519(n595,n583,n594);
not gate_520(n596,n595);
and gate_521(n597,n109,n596);
not gate_522(n598,n597);
and gate_523(n599,n329,n557);
not gate_524(n600,n599);
and gate_525(n601,pi34,n599);
not gate_526(n602,n601);
and gate_527(n603,n598,n602);
not gate_528(n604,n603);
and gate_529(n605,n108,n604);
not gate_530(n606,n605);
and gate_531(n607,n569,n606);
not gate_532(n608,n607);
and gate_533(n609,n105,n608);
not gate_534(n610,n609);
and gate_535(n611,n83,n610);
not gate_536(n612,n611);
and gate_537(po01,pi33,n612);
and gate_538(n614,pi37,n205);
not gate_539(n615,n614);
and gate_540(n616,n110,n193);
not gate_541(n617,n616);
and gate_542(n618,n615,n617);
not gate_543(n619,n618);
and gate_544(n620,n113,n619);
not gate_545(n621,n620);
and gate_546(n622,n217,n496);
not gate_547(n623,n622);
and gate_548(n624,n184,n623);
not gate_549(n625,n624);
and gate_550(n626,n125,n625);
not gate_551(n627,n626);
and gate_552(n628,n621,n627);
not gate_553(n629,n628);
and gate_554(n630,pi34,n629);
not gate_555(n631,n630);
and gate_556(n632,n159,n496);
not gate_557(n633,n632);
and gate_558(n634,n107,n219);
not gate_559(n635,n634);
and gate_560(n636,n633,n635);
not gate_561(n637,n636);
and gate_562(n638,n101,pi30);
not gate_563(n639,n638);
and gate_564(n640,pi29,n639);
not gate_565(n641,n640);
and gate_566(n642,pi28,n103);
not gate_567(n643,n642);
and gate_568(n644,n102,n643);
not gate_569(n645,n644);
and gate_570(n646,n641,n645);
not gate_571(n647,n646);
and gate_572(n648,n637,n647);
not gate_573(n649,n648);
and gate_574(n650,n188,n450);
not gate_575(n651,n650);
and gate_576(n652,n443,n651);
and gate_577(n653,pi15,n652);
and gate_578(n654,pi11,n86);
not gate_579(n655,n654);
and gate_580(n656,n539,n655);
not gate_581(n657,n656);
and gate_582(n658,n107,n657);
and gate_583(n659,n653,n658);
not gate_584(n660,n659);
and gate_585(n661,n649,n660);
not gate_586(n662,n661);
and gate_587(n663,n104,n662);
and gate_588(n664,n81,n663);
not gate_589(n665,n664);
and gate_590(n666,n631,n665);
not gate_591(n667,n666);
and gate_592(n668,n108,n667);
not gate_593(n669,n668);
and gate_594(n670,n200,n487);
not gate_595(n671,n670);
and gate_596(n672,n275,n671);
not gate_597(n673,n672);
and gate_598(n674,pi09,n359);
not gate_599(n675,n674);
and gate_600(n676,n355,n675);
not gate_601(n677,n676);
and gate_602(n678,n196,n677);
and gate_603(n679,pi24,n678);
and gate_604(n680,pi23,n679);
and gate_605(n681,n341,n680);
and gate_606(n682,pi15,n681);
not gate_607(n683,n682);
and gate_608(n684,n496,n682);
not gate_609(n685,n684);
and gate_610(n686,n673,n685);
not gate_611(n687,n686);
and gate_612(n688,n112,n687);
not gate_613(n689,n688);
and gate_614(n690,pi40,n340);
not gate_615(n691,n690);
and gate_616(n692,pi22,n485);
and gate_617(n693,n690,n692);
and gate_618(n694,n95,n693);
and gate_619(n695,pi15,n694);
not gate_620(n696,n695);
and gate_621(n697,n181,n695);
not gate_622(n698,n697);
and gate_623(n699,n689,n698);
not gate_624(n700,n699);
and gate_625(n701,n81,n700);
not gate_626(n702,n701);
and gate_627(n703,pi38,n400);
not gate_628(n704,n703);
and gate_629(n705,n330,n704);
not gate_630(n706,n705);
and gate_631(n707,pi37,n706);
not gate_632(n708,n707);
and gate_633(n709,n702,n708);
not gate_634(n710,n709);
and gate_635(n711,n379,n710);
not gate_636(n712,n711);
and gate_637(n713,n669,n712);
not gate_638(n714,n713);
and gate_639(n715,n109,n714);
not gate_640(n716,n715);
and gate_641(n717,pi37,n468);
not gate_642(n718,n717);
and gate_643(n719,pi38,n414);
not gate_644(n720,n719);
and gate_645(n721,n110,n719);
not gate_646(n722,n721);
and gate_647(n723,n718,n722);
not gate_648(n724,n723);
and gate_649(n725,n108,n724);
not gate_650(n726,n725);
and gate_651(n727,pi35,n159);
not gate_652(n728,n727);
and gate_653(n729,n218,n728);
not gate_654(n730,n729);
and gate_655(n731,pi38,n730);
not gate_656(n732,n731);
and gate_657(n733,pi35,n185);
and gate_658(n734,n388,n733);
not gate_659(n735,n734);
and gate_660(n736,n732,n735);
not gate_661(n737,n736);
and gate_662(n738,n110,n737);
not gate_663(n739,n738);
and gate_664(n740,n726,n739);
not gate_665(n741,n740);
and gate_666(n742,pi36,n741);
not gate_667(n743,n742);
and gate_668(n744,n219,n547);
not gate_669(n745,n744);
and gate_670(n746,n743,n745);
not gate_671(n747,n746);
and gate_672(n748,n107,n747);
not gate_673(n749,n748);
and gate_674(n750,n716,n749);
not gate_675(n751,n750);
and gate_676(n752,n105,n751);
not gate_677(n753,n752);
and gate_678(n754,n83,n753);
not gate_679(n755,n754);
and gate_680(po02,pi33,n755);
and gate_681(n757,pi21,pi22);
not gate_682(n758,n757);
and gate_683(n759,n196,n758);
and gate_684(n760,pi15,n759);
and gate_685(n761,n81,n760);
not gate_686(n762,n761);
and gate_687(n763,pi39,n762);
not gate_688(n764,n763);
and gate_689(n765,pi40,n764);
not gate_690(n766,n765);
and gate_691(n767,n112,n126);
not gate_692(n768,n767);
and gate_693(n769,n766,n768);
not gate_694(n770,n769);
and gate_695(n771,n496,n770);
not gate_696(n772,n771);
and gate_697(n773,n218,n447);
not gate_698(n774,n773);
and gate_699(n775,n772,n774);
and gate_700(n776,n80,n110);
and gate_701(n777,n327,n776);
not gate_702(n778,n777);
and gate_703(n779,n110,n113);
not gate_704(n780,n779);
and gate_705(n781,n186,n780);
not gate_706(n782,n781);
and gate_707(n783,pi02,n143);
not gate_708(n784,n783);
and gate_709(n785,n782,n783);
not gate_710(n786,n785);
and gate_711(n787,n778,n786);
not gate_712(n788,n787);
and gate_713(n789,pi00,n77);
and gate_714(n790,n788,n789);
not gate_715(n791,n790);
and gate_716(n792,n775,n791);
not gate_717(n793,n792);
and gate_718(n794,pi34,n793);
not gate_719(n795,n794);
and gate_720(n796,pi40,n262);
not gate_721(n797,n796);
and gate_722(n798,pi11,n797);
not gate_723(n799,n798);
and gate_724(n800,n81,n799);
not gate_725(n801,n800);
and gate_726(n802,n263,n432);
not gate_727(n803,n802);
and gate_728(n804,pi40,n802);
not gate_729(n805,n804);
and gate_730(n806,n455,n804);
not gate_731(n807,n806);
and gate_732(n808,n801,n807);
not gate_733(n809,n808);
and gate_734(n810,n110,n809);
not gate_735(n811,n810);
and gate_736(n812,n88,pi17);
and gate_737(n813,pi11,n812);
not gate_738(n814,n813);
and gate_739(n815,n107,n814);
and gate_740(n816,n84,n815);
and gate_741(n817,n81,n816);
not gate_742(n818,n817);
and gate_743(n819,n811,n818);
not gate_744(n820,n819);
and gate_745(n821,pi39,n820);
not gate_746(n822,n821);
and gate_747(n823,n81,n254);
and gate_748(n824,n110,n327);
not gate_749(n825,n824);
and gate_750(n826,n823,n824);
not gate_751(n827,n826);
and gate_752(n828,n822,n827);
not gate_753(n829,n828);
and gate_754(n830,pi38,n829);
not gate_755(n831,n830);
and gate_756(n832,n91,n112);
not gate_757(n833,n832);
and gate_758(n834,pi16,n833);
not gate_759(n835,n834);
and gate_760(n836,n84,n835);
not gate_761(n837,n836);
and gate_762(n838,pi11,n263);
not gate_763(n839,n838);
and gate_764(n840,n112,n839);
not gate_765(n841,n840);
and gate_766(n842,n837,n841);
not gate_767(n843,n842);
and gate_768(n844,pi37,n843);
not gate_769(n845,n844);
and gate_770(n846,n90,pi40);
and gate_771(n847,n84,n846);
not gate_772(n848,n847);
and gate_773(n849,n845,n848);
not gate_774(n850,n849);
and gate_775(n851,n111,n850);
not gate_776(n852,n851);
and gate_777(n853,pi39,n254);
not gate_778(n854,n853);
and gate_779(n855,n852,n854);
not gate_780(n856,n855);
and gate_781(n857,n107,n856);
and gate_782(n858,n81,n857);
not gate_783(n859,n858);
and gate_784(n860,n831,n859);
not gate_785(n861,n860);
and gate_786(n862,pi12,n861);
not gate_787(n863,n862);
and gate_788(n864,n185,n221);
not gate_789(n865,n864);
and gate_790(n866,n184,n865);
not gate_791(n867,n866);
and gate_792(n868,n86,n867);
not gate_793(n869,n868);
and gate_794(n870,n107,n468);
not gate_795(n871,n870);
and gate_796(n872,n573,n871);
not gate_797(n873,n872);
and gate_798(n874,n254,n873);
not gate_799(n875,n874);
and gate_800(n876,n869,n875);
not gate_801(n877,n876);
and gate_802(n878,pi11,n877);
not gate_803(n879,n878);
and gate_804(n880,n159,n447);
not gate_805(n881,n880);
and gate_806(n882,n86,n880);
not gate_807(n883,n882);
and gate_808(n884,n879,n883);
not gate_809(n885,n884);
and gate_810(n886,n81,n885);
not gate_811(n887,n886);
and gate_812(n888,n863,n887);
not gate_813(n889,n888);
and gate_814(n890,pi15,n889);
not gate_815(n891,n890);
and gate_816(n892,n86,pi15);
not gate_817(n893,n892);
and gate_818(n894,n159,n893);
and gate_819(n895,n84,n894);
not gate_820(n896,n895);
and gate_821(n897,n101,n231);
not gate_822(n898,n897);
and gate_823(n899,n217,n898);
not gate_824(n900,n899);
and gate_825(n901,n104,n900);
and gate_826(n902,n896,n901);
not gate_827(n903,n902);
and gate_828(n904,pi38,n903);
not gate_829(n905,n904);
and gate_830(n906,pi12,pi14);
and gate_831(n907,pi15,n130);
and gate_832(n908,n906,n907);
not gate_833(n909,n908);
and gate_834(n910,pi31,n909);
not gate_835(n911,n910);
and gate_836(n912,n905,n911);
not gate_837(n913,n912);
and gate_838(n914,n107,n913);
not gate_839(n915,n914);
and gate_840(n916,n623,n881);
not gate_841(n917,n916);
and gate_842(n918,n89,n917);
not gate_843(n919,n918);
and gate_844(n920,n373,n444);
not gate_845(n921,n920);
and gate_846(n922,n919,n921);
not gate_847(n923,n922);
and gate_848(n924,n87,n923);
not gate_849(n925,n924);
and gate_850(n926,n915,n925);
not gate_851(n927,n926);
and gate_852(n928,n81,n927);
not gate_853(n929,n928);
and gate_854(n930,n891,n929);
and gate_855(n931,n795,n930);
not gate_856(n932,n931);
and gate_857(n933,n108,n932);
not gate_858(n934,n933);
and gate_859(n935,n184,n186);
not gate_860(n936,n935);
and gate_861(n937,n98,n936);
not gate_862(n938,n937);
and gate_863(n939,n110,n328);
not gate_864(n940,n939);
and gate_865(n941,n758,n940);
and gate_866(n942,n111,n941);
not gate_867(n943,n942);
and gate_868(n944,n92,n95);
and gate_869(n945,n84,n944);
not gate_870(n946,n945);
and gate_871(n947,pi22,n946);
not gate_872(n948,n947);
and gate_873(n949,n183,n948);
not gate_874(n950,n949);
and gate_875(n951,n943,n950);
and gate_876(n952,n938,n951);
not gate_877(n953,n952);
and gate_878(n954,n197,n953);
and gate_879(n955,n81,n954);
not gate_880(n956,n955);
and gate_881(n957,n111,n218);
not gate_882(n958,n957);
and gate_883(n959,pi00,n159);
not gate_884(n960,n959);
and gate_885(n961,n958,n960);
not gate_886(n962,n961);
and gate_887(n963,pi37,n962);
not gate_888(n964,n963);
and gate_889(n965,n956,n964);
not gate_890(n966,n965);
and gate_891(n967,n379,n966);
not gate_892(n968,n967);
and gate_893(n969,n934,n968);
not gate_894(n970,n969);
and gate_895(n971,n109,n970);
not gate_896(n972,n971);
and gate_897(n973,n110,n182);
not gate_898(n974,n973);
and gate_899(n975,n126,n974);
and gate_900(n976,pi00,n975);
not gate_901(n977,n976);
and gate_902(n978,pi39,n538);
not gate_903(n979,n978);
and gate_904(n980,n110,n979);
not gate_905(n981,n980);
and gate_906(n982,n111,n981);
not gate_907(n983,n982);
and gate_908(n984,n977,n983);
not gate_909(n985,n984);
and gate_910(n986,pi40,n985);
not gate_911(n987,n986);
and gate_912(n988,pi37,pi39);
not gate_913(n989,n988);
and gate_914(n990,n110,n526);
and gate_915(n991,n412,n990);
not gate_916(n992,n991);
and gate_917(n993,n989,n992);
and gate_918(n994,n987,n993);
not gate_919(n995,n994);
and gate_920(n996,n108,n995);
not gate_921(n997,n996);
and gate_922(n998,pi35,n327);
not gate_923(n999,n998);
and gate_924(n1000,n704,n999);
not gate_925(n1001,n1000);
and gate_926(n1002,n80,n1001);
not gate_927(n1003,n1002);
and gate_928(n1004,pi04,pi38);
and gate_929(n1005,n114,n1004);
not gate_930(n1006,n1005);
and gate_931(n1007,pi35,n1005);
not gate_932(n1008,n1007);
and gate_933(n1009,n1003,n1008);
not gate_934(n1010,n1009);
and gate_935(n1011,pi37,n1010);
and gate_936(n1012,n789,n1011);
not gate_937(n1013,n1012);
and gate_938(n1014,n160,n218);
not gate_939(n1015,n1014);
and gate_940(n1016,pi38,n1015);
not gate_941(n1017,n1016);
and gate_942(n1018,n99,n185);
not gate_943(n1019,n1018);
and gate_944(n1020,n1017,n1019);
not gate_945(n1021,n1020);
and gate_946(n1022,n547,n1021);
not gate_947(n1023,n1022);
and gate_948(n1024,n1013,n1023);
and gate_949(n1025,n997,n1024);
not gate_950(n1026,n1025);
and gate_951(n1027,pi36,n1026);
not gate_952(n1028,n1027);
and gate_953(n1029,pi21,pi23);
not gate_954(n1030,n1029);
and gate_955(n1031,n447,n1030);
and gate_956(n1032,n197,n1031);
and gate_957(n1033,n81,n1032);
not gate_958(n1034,n1033);
and gate_959(n1035,n497,n1034);
not gate_960(n1036,n1035);
and gate_961(n1037,pi39,n1036);
not gate_962(n1038,n1037);
and gate_963(n1039,pi37,n146);
and gate_964(n1040,pi00,n1039);
not gate_965(n1041,n1040);
and gate_966(n1042,n1038,n1041);
not gate_967(n1043,n1042);
and gate_968(n1044,pi35,n1043);
not gate_969(n1045,n1044);
and gate_970(n1046,n81,pi37);
and gate_971(n1047,n205,n1046);
not gate_972(n1048,n1047);
and gate_973(n1049,n1045,n1048);
not gate_974(n1050,n1049);
and gate_975(n1051,n113,n1050);
not gate_976(n1052,n1051);
and gate_977(n1053,n84,n108);
and gate_978(n1054,n181,n1053);
and gate_979(n1055,n1046,n1054);
not gate_980(n1056,n1055);
and gate_981(n1057,n1052,n1056);
and gate_982(n1058,n1028,n1057);
not gate_983(n1059,n1058);
and gate_984(n1060,n107,n1059);
not gate_985(n1061,n1060);
and gate_986(n1062,n972,n1061);
not gate_987(n1063,n1062);
and gate_988(n1064,n105,n1063);
not gate_989(n1065,n1064);
and gate_990(n1066,n83,n1065);
not gate_991(n1067,n1066);
and gate_992(po03,pi33,n1067);
and gate_993(n1069,n109,n147);
not gate_994(n1070,n1069);
and gate_995(n1071,pi36,n217);
not gate_996(n1072,n1071);
and gate_997(n1073,n394,n1072);
not gate_998(n1074,n1073);
and gate_999(n1075,n77,n80);
not gate_1000(n1076,n1075);
and gate_1001(n1077,n1074,n1075);
not gate_1002(n1078,n1077);
and gate_1003(n1079,n1070,n1078);
not gate_1004(n1080,n1079);
and gate_1005(n1081,pi00,n1080);
not gate_1006(n1082,n1081);
and gate_1007(n1083,pi36,pi40);
not gate_1008(n1084,n1083);
and gate_1009(n1085,pi39,n1084);
and gate_1010(n1086,n297,n696);
not gate_1011(n1087,n1086);
and gate_1012(n1088,n81,n1087);
not gate_1013(n1089,n1088);
and gate_1014(n1090,n109,n1089);
not gate_1015(n1091,n1090);
and gate_1016(n1092,n1085,n1091);
and gate_1017(n1093,n110,n1092);
not gate_1018(n1094,n1093);
and gate_1019(n1095,n1082,n1094);
not gate_1020(n1096,n1095);
and gate_1021(n1097,pi38,n1096);
not gate_1022(n1098,n1097);
and gate_1023(n1099,n297,n683);
not gate_1024(n1100,n1099);
and gate_1025(n1101,n81,n1100);
not gate_1026(n1102,n1101);
and gate_1027(n1103,n112,n1102);
not gate_1028(n1104,n1103);
and gate_1029(n1105,pi37,pi40);
not gate_1030(n1106,n1105);
and gate_1031(n1107,n1104,n1105);
and gate_1032(n1108,n109,n1107);
not gate_1033(n1109,n1108);
and gate_1034(n1110,n297,n495);
and gate_1035(n1111,n336,n1110);
not gate_1036(n1112,n1111);
and gate_1037(n1113,n109,n1112);
and gate_1038(n1114,n81,n1113);
not gate_1039(n1115,n1114);
and gate_1040(n1116,n99,pi26);
not gate_1041(n1117,n1116);
and gate_1042(n1118,pi36,n1117);
not gate_1043(n1119,n1118);
and gate_1044(n1120,n1115,n1119);
not gate_1045(n1121,n1120);
and gate_1046(n1122,n389,n1121);
not gate_1047(n1123,n1122);
and gate_1048(n1124,n1109,n1123);
not gate_1049(n1125,n1124);
and gate_1050(n1126,n111,n1125);
not gate_1051(n1127,n1126);
and gate_1052(n1128,n156,n327);
not gate_1053(n1129,n1128);
and gate_1054(n1130,n1127,n1129);
and gate_1055(n1131,n1098,n1130);
not gate_1056(n1132,n1131);
and gate_1057(n1133,pi35,n1132);
not gate_1058(n1134,n1133);
and gate_1059(n1135,n111,n131);
not gate_1060(n1136,n1135);
and gate_1061(n1137,pi38,n403);
not gate_1062(n1138,n1137);
and gate_1063(n1139,n434,n1138);
and gate_1064(n1140,n1136,n1139);
and gate_1065(n1141,n432,n1140);
not gate_1066(n1142,n1141);
and gate_1067(n1143,pi31,n1142);
not gate_1068(n1144,n1143);
and gate_1069(n1145,pi11,n906);
not gate_1070(n1146,n1145);
and gate_1071(n1147,n196,n443);
and gate_1072(n1148,n1146,n1147);
and gate_1073(n1149,pi38,n1148);
and gate_1074(n1150,pi15,n1149);
not gate_1075(n1151,n1150);
and gate_1076(n1152,n111,n199);
not gate_1077(n1153,n1152);
and gate_1078(n1154,n1151,n1153);
not gate_1079(n1155,n1154);
and gate_1080(n1156,n128,n1155);
not gate_1081(n1157,n1156);
and gate_1082(n1158,n193,n897);
not gate_1083(n1159,n1158);
and gate_1084(n1160,n1157,n1159);
not gate_1085(n1161,n1160);
and gate_1086(n1162,pi40,n1161);
not gate_1087(n1163,n1162);
and gate_1088(n1164,n187,n1148);
and gate_1089(n1165,pi15,n1164);
not gate_1090(n1166,n1165);
and gate_1091(n1167,n1163,n1166);
and gate_1092(n1168,n1144,n1167);
not gate_1093(n1169,n1168);
and gate_1094(n1170,n109,n1169);
and gate_1095(n1171,n81,n1170);
not gate_1096(n1172,n1171);
and gate_1097(n1173,n111,pi40);
not gate_1098(n1174,n1173);
and gate_1099(n1175,n411,n1174);
not gate_1100(n1176,n1175);
and gate_1101(n1177,pi37,n1176);
not gate_1102(n1178,n1177);
and gate_1103(n1179,n538,n1173);
not gate_1104(n1180,n1179);
and gate_1105(n1181,n1178,n1180);
not gate_1106(n1182,n1181);
and gate_1107(n1183,pi39,n1182);
not gate_1108(n1184,n1183);
and gate_1109(n1185,n722,n1184);
not gate_1110(n1186,n1185);
and gate_1111(n1187,pi36,n1186);
not gate_1112(n1188,n1187);
and gate_1113(n1189,n1172,n1188);
not gate_1114(n1190,n1189);
and gate_1115(n1191,n108,n1190);
not gate_1116(n1192,n1191);
and gate_1117(n1193,n219,n557);
not gate_1118(n1194,n1193);
and gate_1119(n1195,n1192,n1194);
and gate_1120(n1196,n1134,n1195);
not gate_1121(n1197,n1196);
and gate_1122(n1198,n107,n1197);
not gate_1123(n1199,n1198);
and gate_1124(n1200,n80,n328);
not gate_1125(n1201,n1200);
and gate_1126(n1202,pi40,n390);
not gate_1127(n1203,n1202);
and gate_1128(n1204,n1200,n1203);
and gate_1129(n1205,n789,n1204);
not gate_1130(n1206,n1205);
and gate_1131(n1207,n81,n296);
not gate_1132(n1208,n1207);
and gate_1133(n1209,pi40,n1208);
not gate_1134(n1210,n1209);
and gate_1135(n1211,n988,n1210);
not gate_1136(n1212,n1211);
and gate_1137(n1213,n1206,n1212);
not gate_1138(n1214,n1213);
and gate_1139(n1215,pi34,n1214);
not gate_1140(n1216,n1215);
and gate_1141(n1217,n393,n647);
and gate_1142(n1218,n81,n1217);
not gate_1143(n1219,n1218);
and gate_1144(n1220,n1216,n1219);
not gate_1145(n1221,n1220);
and gate_1146(n1222,n111,n1221);
not gate_1147(n1223,n1222);
and gate_1148(n1224,pi34,n990);
not gate_1149(n1225,n1224);
and gate_1150(n1226,n1223,n1225);
not gate_1151(n1227,n1226);
and gate_1152(n1228,n109,n1227);
not gate_1153(n1229,n1228);
and gate_1154(n1230,n602,n1229);
not gate_1155(n1231,n1230);
and gate_1156(n1232,n108,n1231);
not gate_1157(n1233,n1232);
and gate_1158(n1234,n1199,n1233);
not gate_1159(n1235,n1234);
and gate_1160(po04,n429,n1235);
and gate_1161(n1237,n96,n379);
and gate_1162(n1238,n197,n1237);
and gate_1163(n1239,n81,n1238);
not gate_1164(n1240,n1239);
and gate_1165(n1241,pi34,n127);
not gate_1166(n1242,n1241);
and gate_1167(n1243,n1240,n1242);
not gate_1168(n1244,n1243);
and gate_1169(n1245,n190,n1244);
not gate_1170(n1246,n1245);
and gate_1171(n1247,pi40,n758);
and gate_1172(n1248,n264,n1247);
and gate_1173(n1249,pi15,n1248);
and gate_1174(n1250,n81,n1249);
not gate_1175(n1251,n1250);
and gate_1176(n1252,n80,n113);
not gate_1177(n1253,n1252);
and gate_1178(n1254,n114,n1253);
not gate_1179(n1255,n1254);
and gate_1180(n1256,n1201,n1255);
not gate_1181(n1257,n1256);
and gate_1182(n1258,n110,n1257);
and gate_1183(n1259,n789,n1258);
not gate_1184(n1260,n1259);
and gate_1185(n1261,n1251,n1260);
not gate_1186(n1262,n1261);
and gate_1187(n1263,pi34,n1262);
not gate_1188(n1264,n1263);
and gate_1189(n1265,pi13,n291);
not gate_1190(n1266,n1265);
and gate_1191(n1267,n107,n1265);
not gate_1192(n1268,n1267);
and gate_1193(n1269,n403,n1268);
not gate_1194(n1270,n1269);
and gate_1195(n1271,n198,n1270);
not gate_1196(n1272,n1271);
and gate_1197(n1273,n130,n803);
not gate_1198(n1274,n1273);
and gate_1199(n1275,n848,n1274);
not gate_1200(n1276,n1275);
and gate_1201(n1277,n196,n1276);
not gate_1202(n1278,n1277);
and gate_1203(n1279,pi12,n88);
and gate_1204(n1280,pi11,n1279);
and gate_1205(n1281,n130,n1280);
not gate_1206(n1282,n1281);
and gate_1207(n1283,n1278,n1282);
not gate_1208(n1284,n1283);
and gate_1209(n1285,n107,n1284);
and gate_1210(n1286,pi15,n1285);
not gate_1211(n1287,n1286);
and gate_1212(n1288,n1272,n1287);
not gate_1213(n1289,n1288);
and gate_1214(n1290,n104,n1289);
and gate_1215(n1291,n81,n1290);
not gate_1216(n1292,n1291);
and gate_1217(n1293,n1264,n1292);
not gate_1218(n1294,n1293);
and gate_1219(n1295,n111,n1294);
not gate_1220(n1296,n1295);
and gate_1221(n1297,n107,pi39);
not gate_1222(n1298,n1297);
and gate_1223(n1299,n527,n1298);
not gate_1224(n1300,n1299);
and gate_1225(n1301,n84,n1300);
not gate_1226(n1302,n1301);
and gate_1227(n1303,pi38,pi40);
not gate_1228(n1304,n1303);
and gate_1229(n1305,n91,pi39);
not gate_1230(n1306,n1305);
and gate_1231(n1307,n1303,n1305);
not gate_1232(n1308,n1307);
and gate_1233(n1309,n1302,n1308);
not gate_1234(n1310,n1309);
and gate_1235(n1311,n196,n1310);
and gate_1236(n1312,n90,n1311);
not gate_1237(n1313,n1312);
and gate_1238(n1314,n703,n1280);
not gate_1239(n1315,n1314);
and gate_1240(n1316,n1313,n1315);
not gate_1241(n1317,n1316);
and gate_1242(n1318,pi15,n1317);
not gate_1243(n1319,n1318);
and gate_1244(n1320,pi11,n245);
not gate_1245(n1321,n1320);
and gate_1246(n1322,n161,n1321);
and gate_1247(n1323,n107,n1322);
not gate_1248(n1324,n1323);
and gate_1249(n1325,n296,n1300);
not gate_1250(n1326,n1325);
and gate_1251(n1327,n1324,n1326);
and gate_1252(n1328,n1319,n1327);
not gate_1253(n1329,n1328);
and gate_1254(n1330,n104,n1329);
and gate_1255(n1331,n81,n1330);
not gate_1256(n1332,n1331);
and gate_1257(n1333,n401,n527);
not gate_1258(n1334,n1333);
and gate_1259(n1335,pi34,n1334);
not gate_1260(n1336,n1335);
and gate_1261(n1337,n1332,n1336);
not gate_1262(n1338,n1337);
and gate_1263(n1339,n110,n1338);
not gate_1264(n1340,n1339);
and gate_1265(n1341,n230,n232);
not gate_1266(n1342,n1341);
and gate_1267(n1343,n217,n1342);
not gate_1268(n1344,n1343);
and gate_1269(n1345,n285,n1344);
not gate_1270(n1346,n1345);
and gate_1271(n1347,pi38,n1346);
and gate_1272(n1348,n107,n1347);
and gate_1273(n1349,n104,n1348);
and gate_1274(n1350,n81,n1349);
not gate_1275(n1351,n1350);
and gate_1276(n1352,n1340,n1351);
and gate_1277(n1353,n1296,n1352);
not gate_1278(n1354,n1353);
and gate_1279(n1355,n108,n1354);
not gate_1280(n1356,n1355);
and gate_1281(n1357,pi21,pi24);
not gate_1282(n1358,n1357);
and gate_1283(n1359,n264,n1358);
and gate_1284(n1360,n447,n1359);
and gate_1285(n1361,pi15,n1360);
not gate_1286(n1362,n1361);
and gate_1287(n1363,n87,n110);
not gate_1288(n1364,n1363);
and gate_1289(n1365,n494,n1363);
not gate_1290(n1366,n1365);
and gate_1291(n1367,pi37,n362);
not gate_1292(n1368,n1367);
and gate_1293(n1369,pi40,n1368);
not gate_1294(n1370,n1369);
and gate_1295(n1371,n95,n1370);
not gate_1296(n1372,n1371);
and gate_1297(n1373,n96,n113);
not gate_1298(n1374,n1373);
and gate_1299(n1375,pi24,n1374);
and gate_1300(n1376,n1372,n1375);
not gate_1301(n1377,n1376);
and gate_1302(n1378,n197,n1377);
not gate_1303(n1379,n1378);
and gate_1304(n1380,n1366,n1379);
not gate_1305(n1381,n1380);
and gate_1306(n1382,n185,n1381);
not gate_1307(n1383,n1382);
and gate_1308(n1384,n1362,n1383);
not gate_1309(n1385,n1384);
and gate_1310(n1386,n81,n1385);
not gate_1311(n1387,n1386);
and gate_1312(n1388,pi00,pi39);
not gate_1313(n1389,n1388);
and gate_1314(n1390,pi38,n1389);
not gate_1315(n1391,n1390);
and gate_1316(n1392,n147,n1391);
not gate_1317(n1393,n1392);
and gate_1318(n1394,n1387,n1393);
not gate_1319(n1395,n1394);
and gate_1320(n1396,n379,n1395);
not gate_1321(n1397,n1396);
and gate_1322(n1398,n1356,n1397);
and gate_1323(n1399,n1246,n1398);
not gate_1324(n1400,n1399);
and gate_1325(n1401,n109,n1400);
not gate_1326(n1402,n1401);
and gate_1327(n1403,n108,pi36);
and gate_1328(n1404,n1303,n1403);
not gate_1329(n1405,n1404);
and gate_1330(n1406,n111,n113);
not gate_1331(n1407,n1406);
and gate_1332(n1408,n118,n1406);
not gate_1333(n1409,n1408);
and gate_1334(n1410,n1405,n1409);
not gate_1335(n1411,n1410);
and gate_1336(n1412,n585,n1411);
not gate_1337(n1413,n1412);
and gate_1338(n1414,pi01,pi04);
not gate_1339(n1415,n1414);
and gate_1340(n1416,n194,n1415);
and gate_1341(n1417,pi38,n1076);
not gate_1342(n1418,n1417);
and gate_1343(n1419,n1416,n1418);
and gate_1344(n1420,n147,n1419);
and gate_1345(n1421,pi35,n1420);
not gate_1346(n1422,n1421);
and gate_1347(n1423,n80,n217);
not gate_1348(n1424,n1423);
and gate_1349(n1425,n784,n1424);
not gate_1350(n1426,n1425);
and gate_1351(n1427,n118,n1426);
and gate_1352(n1428,n77,n1427);
not gate_1353(n1429,n1428);
and gate_1354(n1430,pi40,n1076);
and gate_1355(n1431,n108,n1430);
not gate_1356(n1432,n1431);
and gate_1357(n1433,n1429,n1432);
not gate_1358(n1434,n1433);
and gate_1359(n1435,pi36,pi38);
and gate_1360(n1436,n1434,n1435);
not gate_1361(n1437,n1436);
and gate_1362(n1438,n1422,n1437);
and gate_1363(n1439,n1413,n1438);
not gate_1364(n1440,n1439);
and gate_1365(n1441,pi00,n1440);
not gate_1366(n1442,n1441);
and gate_1367(n1443,pi36,n1173);
not gate_1368(n1444,n1443);
and gate_1369(n1445,pi15,n97);
and gate_1370(n1446,n81,n1445);
and gate_1371(n1447,pi35,n410);
and gate_1372(n1448,n1446,n1447);
not gate_1373(n1449,n1448);
and gate_1374(n1450,n1444,n1449);
not gate_1375(n1451,n1450);
and gate_1376(n1452,n196,n1451);
not gate_1377(n1453,n1452);
and gate_1378(n1454,pi35,pi36);
and gate_1379(n1455,n1304,n1454);
not gate_1380(n1456,n1455);
and gate_1381(n1457,n1453,n1456);
not gate_1382(n1458,n1457);
and gate_1383(n1459,n110,n1458);
not gate_1384(n1460,n1459);
and gate_1385(n1461,pi35,pi40);
not gate_1386(n1462,n1461);
and gate_1387(n1463,pi36,n1175);
and gate_1388(n1464,n1462,n1463);
not gate_1389(n1465,n1464);
and gate_1390(n1466,n104,n898);
and gate_1391(n1467,n81,n1466);
not gate_1392(n1468,n1467);
and gate_1393(n1469,n108,n1468);
not gate_1394(n1470,n1469);
and gate_1395(n1471,n1406,n1470);
not gate_1396(n1472,n1471);
and gate_1397(n1473,n1465,n1472);
not gate_1398(n1474,n1473);
and gate_1399(n1475,pi37,n1474);
not gate_1400(n1476,n1475);
and gate_1401(n1477,n1460,n1476);
not gate_1402(n1478,n1477);
and gate_1403(n1479,pi39,n1478);
not gate_1404(n1480,n1479);
and gate_1405(n1481,n111,n1117);
and gate_1406(n1482,pi35,n1481);
not gate_1407(n1483,n1482);
and gate_1408(n1484,n113,n413);
not gate_1409(n1485,n1484);
and gate_1410(n1486,n193,n1485);
and gate_1411(n1487,n108,n1486);
not gate_1412(n1488,n1487);
and gate_1413(n1489,n1483,n1488);
not gate_1414(n1490,n1489);
and gate_1415(n1491,n110,n1490);
not gate_1416(n1492,n1491);
and gate_1417(n1493,n108,pi37);
not gate_1418(n1494,n1493);
and gate_1419(n1495,n373,n1493);
not gate_1420(n1496,n1495);
and gate_1421(n1497,n1492,n1496);
not gate_1422(n1498,n1497);
and gate_1423(n1499,pi36,n1498);
not gate_1424(n1500,n1499);
and gate_1425(n1501,n1480,n1500);
and gate_1426(n1502,n1442,n1501);
not gate_1427(n1503,n1502);
and gate_1428(n1504,n107,n1503);
not gate_1429(n1505,n1504);
and gate_1430(n1506,n1402,n1505);
not gate_1431(n1507,n1506);
and gate_1432(po05,n429,n1507);
and gate_1433(n1509,n109,pi38);
not gate_1434(n1510,n1509);
and gate_1435(n1511,n217,n1509);
not gate_1436(n1512,n1511);
and gate_1437(n1513,n633,n1512);
not gate_1438(n1514,n1513);
and gate_1439(n1515,n647,n1514);
not gate_1440(n1516,n1515);
and gate_1441(n1517,pi13,n411);
not gate_1442(n1518,n1517);
and gate_1443(n1519,n1174,n1518);
not gate_1444(n1520,n1519);
and gate_1445(n1521,pi39,n1520);
not gate_1446(n1522,n1521);
and gate_1447(n1523,pi13,n526);
not gate_1448(n1524,n1523);
and gate_1449(n1525,n1522,n1524);
not gate_1450(n1526,n1525);
and gate_1451(n1527,n198,n1526);
not gate_1452(n1528,n1527);
and gate_1453(n1529,pi09,n1322);
not gate_1454(n1530,n1529);
and gate_1455(n1531,n1528,n1530);
not gate_1456(n1532,n1531);
and gate_1457(n1533,n110,n1532);
not gate_1458(n1534,n1533);
and gate_1459(n1535,pi37,n217);
not gate_1460(n1536,n1535);
and gate_1461(n1537,n1266,n1536);
not gate_1462(n1538,n1537);
and gate_1463(n1539,n198,n1538);
and gate_1464(n1540,n111,n1539);
not gate_1465(n1541,n1540);
and gate_1466(n1542,n1534,n1541);
not gate_1467(n1543,n1542);
and gate_1468(n1544,n109,n1543);
not gate_1469(n1545,n1544);
and gate_1470(n1546,n1516,n1545);
not gate_1471(n1547,n1546);
and gate_1472(n1548,n108,n1547);
and gate_1473(n1549,n104,n1548);
not gate_1474(n1550,n1549);
and gate_1475(n1551,pi37,n1173);
not gate_1476(n1552,n1551);
and gate_1477(n1553,n184,n1552);
not gate_1478(n1554,n1553);
and gate_1479(n1555,n109,n1554);
not gate_1480(n1556,n1555);
and gate_1481(n1557,n168,n327);
not gate_1482(n1558,n1557);
and gate_1483(n1559,n1556,n1558);
not gate_1484(n1560,n1559);
and gate_1485(n1561,n87,n1560);
not gate_1486(n1562,n1561);
and gate_1487(n1563,n110,n217);
not gate_1488(n1564,n1563);
and gate_1489(n1565,pi13,n1563);
not gate_1490(n1566,n1565);
and gate_1491(n1567,n1562,n1566);
not gate_1492(n1568,n1567);
and gate_1493(n1569,n198,n1568);
not gate_1494(n1570,n1569);
and gate_1495(n1571,pi19,pi23);
and gate_1496(n1572,n496,n1571);
not gate_1497(n1573,n1572);
and gate_1498(n1574,n448,n1573);
not gate_1499(n1575,n1574);
and gate_1500(n1576,n340,n1575);
not gate_1501(n1577,n1576);
and gate_1502(n1578,n448,n497);
not gate_1503(n1579,n1578);
and gate_1504(n1580,pi21,n1579);
not gate_1505(n1581,n1580);
and gate_1506(n1582,pi18,pi23);
and gate_1507(n1583,pi09,n1582);
and gate_1508(n1584,n496,n1583);
not gate_1509(n1585,n1584);
and gate_1510(n1586,n1581,n1585);
and gate_1511(n1587,n1577,n1586);
not gate_1512(n1588,n1587);
and gate_1513(n1589,pi40,n1588);
not gate_1514(n1590,n1589);
and gate_1515(n1591,n183,n1029);
not gate_1516(n1592,n1591);
and gate_1517(n1593,n1590,n1592);
not gate_1518(n1594,n1593);
and gate_1519(n1595,n109,n1594);
not gate_1520(n1596,n1595);
and gate_1521(n1597,n110,n185);
not gate_1522(n1598,n1597);
and gate_1523(n1599,pi21,n1597);
not gate_1524(n1600,n1599);
and gate_1525(n1601,n1596,n1600);
not gate_1526(n1602,n1601);
and gate_1527(n1603,pi22,n1602);
not gate_1528(n1604,n1603);
and gate_1529(n1605,n1564,n1604);
not gate_1530(n1606,n1605);
and gate_1531(n1607,n486,n1606);
not gate_1532(n1608,n1607);
and gate_1533(n1609,n1570,n1608);
not gate_1534(n1610,n1609);
and gate_1535(n1611,pi35,n1610);
not gate_1536(n1612,n1611);
and gate_1537(n1613,n1550,n1612);
not gate_1538(n1614,n1613);
and gate_1539(n1615,n81,n1614);
not gate_1540(n1616,n1615);
and gate_1541(n1617,pi35,n390);
and gate_1542(n1618,pi00,n1075);
and gate_1543(n1619,n1617,n1618);
not gate_1544(n1620,n1619);
and gate_1545(n1621,n108,n110);
not gate_1546(n1622,n1621);
and gate_1547(n1623,n414,n1621);
not gate_1548(n1624,n1623);
and gate_1549(n1625,n1620,n1624);
not gate_1550(n1626,n1625);
and gate_1551(n1627,pi38,n1626);
not gate_1552(n1628,n1627);
and gate_1553(n1629,n108,n496);
not gate_1554(n1630,n1629);
and gate_1555(n1631,n548,n1630);
not gate_1556(n1632,n1631);
and gate_1557(n1633,pi39,n1632);
not gate_1558(n1634,n1633);
and gate_1559(n1635,n1628,n1634);
not gate_1560(n1636,n1635);
and gate_1561(n1637,n113,n1636);
not gate_1562(n1638,n1637);
and gate_1563(n1639,n219,n1618);
not gate_1564(n1640,n1639);
and gate_1565(n1641,n169,n1640);
not gate_1566(n1642,n1641);
and gate_1567(n1643,pi35,n1642);
not gate_1568(n1644,n1643);
and gate_1569(n1645,pi11,n110);
and gate_1570(n1646,n111,n400);
not gate_1571(n1647,n1646);
and gate_1572(n1648,n1645,n1646);
not gate_1573(n1649,n1648);
and gate_1574(n1650,n1644,n1649);
and gate_1575(n1651,n1638,n1650);
not gate_1576(n1652,n1651);
and gate_1577(n1653,pi36,n1652);
not gate_1578(n1654,n1653);
and gate_1579(n1655,n156,n205);
not gate_1580(n1656,n1655);
and gate_1581(n1657,n217,n447);
not gate_1582(n1658,n1657);
and gate_1583(n1659,n1656,n1658);
not gate_1584(n1660,n1659);
and gate_1585(n1661,pi35,n1660);
not gate_1586(n1662,n1661);
and gate_1587(n1663,n1654,n1662);
and gate_1588(n1664,n1616,n1663);
not gate_1589(n1665,n1664);
and gate_1590(n1666,n107,n1665);
not gate_1591(n1667,n1666);
and gate_1592(n1668,n197,n757);
not gate_1593(n1669,n1668);
and gate_1594(n1670,n200,n1669);
not gate_1595(n1671,n1670);
and gate_1596(n1672,n81,n1671);
not gate_1597(n1673,n1672);
and gate_1598(n1674,n205,n1672);
not gate_1599(n1675,n1674);
and gate_1600(n1676,n194,n1675);
not gate_1601(n1677,n1676);
and gate_1602(n1678,pi37,n1677);
not gate_1603(n1679,n1678);
and gate_1604(n1680,n181,n776);
and gate_1605(n1681,n586,n1680);
not gate_1606(n1682,n1681);
and gate_1607(n1683,n1679,n1682);
not gate_1608(n1684,n1683);
and gate_1609(n1685,pi40,n1684);
and gate_1610(n1686,pi34,n170);
and gate_1611(n1687,n1685,n1686);
not gate_1612(n1688,n1687);
and gate_1613(n1689,n1667,n1688);
not gate_1614(n1690,n1689);
and gate_1615(po06,n429,n1690);
and gate_1616(n1692,n443,n657);
and gate_1617(n1693,n112,n1692);
and gate_1618(n1694,n221,n1693);
and gate_1619(n1695,n104,n1694);
not gate_1620(n1696,n1695);
and gate_1621(n1697,pi40,n196);
and gate_1622(n1698,pi39,n1697);
and gate_1623(n1699,pi34,n1698);
and gate_1624(n1700,n757,n1699);
not gate_1625(n1701,n1700);
and gate_1626(n1702,n1696,n1701);
not gate_1627(n1703,n1702);
and gate_1628(n1704,n111,n1703);
not gate_1629(n1705,n1704);
and gate_1630(n1706,n449,n1692);
and gate_1631(n1707,n107,n1706);
and gate_1632(n1708,n104,n1707);
not gate_1633(n1709,n1708);
and gate_1634(n1710,n1705,n1709);
not gate_1635(n1711,n1710);
and gate_1636(n1712,pi15,n1711);
not gate_1637(n1713,n1712);
and gate_1638(n1714,n104,n897);
and gate_1639(n1715,n227,n1714);
not gate_1640(n1716,n1715);
and gate_1641(n1717,n1713,n1716);
not gate_1642(n1718,n1717);
and gate_1643(n1719,n108,n1718);
not gate_1644(n1720,n1719);
and gate_1645(n1721,n187,n1571);
not gate_1646(n1722,n1721);
and gate_1647(n1723,n184,n1722);
not gate_1648(n1724,n1723);
and gate_1649(n1725,n340,n1724);
not gate_1650(n1726,n1725);
and gate_1651(n1727,pi21,n190);
not gate_1652(n1728,n1727);
and gate_1653(n1729,n187,n1583);
not gate_1654(n1730,n1729);
and gate_1655(n1731,n1728,n1730);
and gate_1656(n1732,n1726,n1731);
not gate_1657(n1733,n1732);
and gate_1658(n1734,pi40,n1733);
not gate_1659(n1735,n1734);
and gate_1660(n1736,pi23,n181);
not gate_1661(n1737,n1736);
and gate_1662(n1738,n330,n1737);
not gate_1663(n1739,n1738);
and gate_1664(n1740,n110,n1739);
and gate_1665(n1741,pi21,n1740);
not gate_1666(n1742,n1741);
and gate_1667(n1743,n1735,n1742);
not gate_1668(n1744,n1743);
and gate_1669(n1745,n379,n1744);
and gate_1670(n1746,n692,n1745);
and gate_1671(n1747,pi15,n1746);
not gate_1672(n1748,n1747);
and gate_1673(n1749,n1720,n1748);
not gate_1674(n1750,n1749);
and gate_1675(n1751,n81,n1750);
not gate_1676(n1752,n1751);
and gate_1677(n1753,n111,n401);
not gate_1678(n1754,n1753);
and gate_1679(n1755,n973,n1754);
not gate_1680(n1756,n1755);
and gate_1681(n1757,n220,n1756);
not gate_1682(n1758,n1757);
and gate_1683(n1759,pi34,n108);
and gate_1684(n1760,n1758,n1759);
not gate_1685(n1761,n1760);
and gate_1686(n1762,n1752,n1761);
not gate_1687(n1763,n1762);
and gate_1688(n1764,n109,n1763);
not gate_1689(n1765,n1764);
and gate_1690(n1766,pi35,n1016);
not gate_1691(n1767,n1766);
and gate_1692(n1768,n85,n509);
and gate_1693(n1769,n1646,n1768);
not gate_1694(n1770,n1769);
and gate_1695(n1771,n1767,n1770);
not gate_1696(n1772,n1771);
and gate_1697(n1773,n557,n1772);
and gate_1698(n1774,n107,n1773);
not gate_1699(n1775,n1774);
and gate_1700(n1776,n1765,n1775);
not gate_1701(n1777,n1776);
and gate_1702(n1778,n105,n1777);
not gate_1703(n1779,n1778);
and gate_1704(n1780,n83,n1779);
not gate_1705(n1781,n1780);
and gate_1706(po07,pi33,n1781);
and gate_1707(n1783,pi34,n109);
and gate_1708(n1784,pi37,n193);
and gate_1709(n1785,n1783,n1784);
not gate_1710(n1786,n1785);
and gate_1711(n1787,n205,n557);
and gate_1712(n1788,n107,n1787);
and gate_1713(n1789,n538,n1788);
not gate_1714(n1790,n1789);
and gate_1715(n1791,n1786,n1790);
not gate_1716(n1792,n1791);
and gate_1717(n1793,pi40,n1792);
and gate_1718(n1794,n108,n1793);
and gate_1719(n1795,n105,n1794);
not gate_1720(n1796,n1795);
and gate_1721(n1797,n83,n1796);
not gate_1722(n1798,n1797);
and gate_1723(po08,pi33,n1798);
and gate_1724(n1800,n108,n1692);
and gate_1725(n1801,n104,n1800);
not gate_1726(n1802,n1801);
and gate_1727(n1803,n651,n1801);
not gate_1728(n1804,n1803);
and gate_1729(n1805,n681,n1461);
and gate_1730(n1806,n187,n1805);
not gate_1731(n1807,n1806);
and gate_1732(n1808,n1804,n1807);
not gate_1733(n1809,n1808);
and gate_1734(n1810,pi15,n1809);
not gate_1735(n1811,n1810);
and gate_1736(n1812,n222,n1493);
and gate_1737(n1813,n1714,n1812);
not gate_1738(n1814,n1813);
and gate_1739(n1815,n1811,n1814);
not gate_1740(n1816,n1815);
and gate_1741(n1817,n109,n1816);
and gate_1742(n1818,n107,n1817);
and gate_1743(n1819,n105,n1818);
and gate_1744(n1820,n81,n1819);
not gate_1745(n1821,n1820);
and gate_1746(n1822,n83,n1821);
not gate_1747(n1823,n1822);
and gate_1748(po09,pi33,n1823);
and gate_1749(n1825,n94,n99);
not gate_1750(n1826,n1825);
and gate_1751(n1827,n97,n113);
not gate_1752(n1828,n1827);
and gate_1753(n1829,n181,n1828);
not gate_1754(n1830,n1829);
and gate_1755(n1831,n330,n1830);
not gate_1756(n1832,n1831);
and gate_1757(n1833,n110,n1832);
not gate_1758(n1834,n1833);
and gate_1759(n1835,n623,n1834);
not gate_1760(n1836,n1835);
and gate_1761(n1837,n379,n1836);
and gate_1762(n1838,pi24,n1837);
not gate_1763(n1839,n1838);
and gate_1764(n1840,n1646,n1759);
not gate_1765(n1841,n1840);
and gate_1766(n1842,n1839,n1841);
not gate_1767(n1843,n1842);
and gate_1768(n1844,n196,n1843);
and gate_1769(n1845,n1826,n1844);
and gate_1770(n1846,n757,n1845);
and gate_1771(n1847,pi15,n1846);
and gate_1772(n1848,n81,n1847);
not gate_1773(n1849,n1848);
and gate_1774(n1850,n1755,n1759);
not gate_1775(n1851,n1850);
and gate_1776(n1852,n1849,n1851);
not gate_1777(n1853,n1852);
and gate_1778(n1854,n109,n1853);
and gate_1779(po10,n429,n1854);
and gate_1780(n1856,n1629,n1693);
and gate_1781(n1857,n104,n1856);
not gate_1782(n1858,n1857);
and gate_1783(n1859,pi35,n340);
and gate_1784(n1860,n692,n1859);
and gate_1785(n1861,n95,n1860);
not gate_1786(n1862,n1861);
and gate_1787(n1863,n1802,n1862);
not gate_1788(n1864,n1863);
and gate_1789(n1865,n449,n1864);
not gate_1790(n1866,n1865);
and gate_1791(n1867,n1858,n1866);
not gate_1792(n1868,n1867);
and gate_1793(n1869,n107,n1868);
and gate_1794(n1870,pi15,n1869);
not gate_1795(n1871,n1870);
and gate_1796(n1872,n108,pi38);
not gate_1797(n1873,n1872);
and gate_1798(n1874,n217,n1872);
and gate_1799(n1875,n1714,n1874);
not gate_1800(n1876,n1875);
and gate_1801(n1877,n1871,n1876);
not gate_1802(n1878,n1877);
and gate_1803(n1879,n81,n1878);
not gate_1804(n1880,n1879);
and gate_1805(n1881,n1761,n1880);
not gate_1806(n1882,n1881);
and gate_1807(n1883,n109,n1882);
and gate_1808(po11,n429,n1883);
and gate_1809(n1885,n76,pi05);
not gate_1810(n1886,n1885);
and gate_1811(n1887,n379,n535);
not gate_1812(n1888,n1887);
and gate_1813(n1889,pi36,n1887);
not gate_1814(n1890,n1889);
and gate_1815(n1891,n109,n110);
not gate_1816(n1892,n1891);
and gate_1817(n1893,n1759,n1891);
not gate_1818(n1894,n1893);
and gate_1819(n1895,n111,n1893);
not gate_1820(n1896,n1895);
and gate_1821(n1897,n1890,n1896);
not gate_1822(n1898,n1897);
and gate_1823(n1899,n113,n1898);
and gate_1824(n1900,pi33,n1899);
and gate_1825(n1901,pi08,n1900);
and gate_1826(n1902,n428,n1901);
and gate_1827(po12,n1885,n1902);
and gate_1828(n1904,n527,n1647);
not gate_1829(n1905,n1904);
and gate_1830(n1906,n109,n1905);
not gate_1831(n1907,n1906);
and gate_1832(n1908,pi36,n185);
not gate_1833(n1909,n1908);
and gate_1834(n1910,n1907,n1909);
not gate_1835(n1911,n1910);
and gate_1836(n1912,n547,n1911);
and gate_1837(n1913,n107,n1912);
and gate_1838(n1914,n105,n1913);
not gate_1839(n1915,n1914);
and gate_1840(n1916,n83,n1915);
not gate_1841(n1917,n1916);
and gate_1842(po13,pi33,n1917);
and gate_1843(n1919,pi13,n1908);
not gate_1844(n1920,n1919);
and gate_1845(n1921,n1907,n1920);
not gate_1846(n1922,n1921);
and gate_1847(n1923,n547,n1922);
and gate_1848(n1924,n107,n1923);
and gate_1849(n1925,n105,n1924);
not gate_1850(n1926,n1925);
and gate_1851(n1927,n83,n1926);
not gate_1852(n1928,n1927);
and gate_1853(po14,pi33,n1928);
and gate_1854(po15,pi07,pi33);
and gate_1855(n1931,n131,n403);
not gate_1856(n1932,n1931);
and gate_1857(n1933,n125,n1932);
and gate_1858(n1934,pi00,n1933);
not gate_1859(n1935,n1934);
and gate_1860(n1936,pi37,n327);
not gate_1861(n1937,n1936);
and gate_1862(n1938,n1935,n1937);
not gate_1863(n1939,n1938);
and gate_1864(n1940,pi38,n1939);
not gate_1865(n1941,n1940);
and gate_1866(n1942,pi40,n195);
not gate_1867(n1943,n1942);
and gate_1868(n1944,pi39,n1943);
not gate_1869(n1945,n1944);
and gate_1870(n1946,n168,n1945);
not gate_1871(n1947,n1946);
and gate_1872(n1948,n1941,n1947);
not gate_1873(n1949,n1948);
and gate_1874(n1950,n108,n1949);
not gate_1875(n1951,n1950);
and gate_1876(n1952,n118,n329);
and gate_1877(n1953,pi00,n142);
and gate_1878(n1954,n143,n1953);
not gate_1879(n1955,n1954);
and gate_1880(n1956,n1952,n1954);
not gate_1881(n1957,n1956);
and gate_1882(n1958,n1951,n1957);
not gate_1883(n1959,n1958);
and gate_1884(n1960,pi36,n1959);
not gate_1885(n1961,n1960);
and gate_1886(n1962,n158,n219);
not gate_1887(n1963,n1962);
and gate_1888(n1964,n1961,n1963);
not gate_1889(n1965,n1964);
and gate_1890(n1966,n107,n1965);
not gate_1891(n1967,n1966);
and gate_1892(n1968,n159,n535);
and gate_1893(n1969,n1686,n1968);
not gate_1894(n1970,n1969);
and gate_1895(n1971,n1967,n1970);
not gate_1896(n1972,n1971);
and gate_1897(po16,n429,n1972);
and gate_1898(n1974,pi39,n780);
not gate_1899(n1975,n1974);
and gate_1900(n1976,n143,n1975);
and gate_1901(n1977,n789,n1976);
not gate_1902(n1978,n1977);
and gate_1903(n1979,n131,n1978);
not gate_1904(n1980,n1979);
and gate_1905(n1981,pi02,n1980);
not gate_1906(n1982,n1981);
and gate_1907(n1983,n77,n124);
not gate_1908(n1984,n1983);
and gate_1909(n1985,n112,n1984);
not gate_1910(n1986,n1985);
and gate_1911(n1987,n1251,n1986);
not gate_1912(n1988,n1987);
and gate_1913(n1989,pi37,n1988);
not gate_1914(n1990,n1989);
and gate_1915(n1991,n1982,n1990);
not gate_1916(n1992,n1991);
and gate_1917(n1993,pi34,n1992);
not gate_1918(n1994,n1993);
and gate_1919(n1995,n159,n236);
not gate_1920(n1996,n1995);
and gate_1921(n1997,n112,n803);
and gate_1922(n1998,n197,n1997);
not gate_1923(n1999,n1998);
and gate_1924(n2000,n1996,n1999);
not gate_1925(n2001,n2000);
and gate_1926(n2002,pi37,n2001);
not gate_1927(n2003,n2002);
and gate_1928(n2004,n197,n847);
not gate_1929(n2005,n2004);
and gate_1930(n2006,n2003,n2005);
not gate_1931(n2007,n2006);
and gate_1932(n2008,n107,n2007);
and gate_1933(n2009,n104,n2008);
and gate_1934(n2010,n81,n2009);
not gate_1935(n2011,n2010);
and gate_1936(n2012,n1994,n2011);
not gate_1937(n2013,n2012);
and gate_1938(n2014,n111,n2013);
not gate_1939(n2015,n2014);
and gate_1940(n2016,n110,n264);
and gate_1941(n2017,n262,n2016);
and gate_1942(n2018,pi15,n2017);
not gate_1943(n2019,n2018);
and gate_1944(n2020,n112,n236);
not gate_1945(n2021,n2020);
and gate_1946(n2022,n2019,n2021);
not gate_1947(n2023,n2022);
and gate_1948(n2024,pi40,n2023);
not gate_1949(n2025,n2024);
and gate_1950(n2026,pi39,n276);
not gate_1951(n2027,n2026);
and gate_1952(n2028,n112,n780);
not gate_1953(n2029,n2028);
and gate_1954(n2030,n90,n2029);
not gate_1955(n2031,n2030);
and gate_1956(n2032,n1306,n2031);
not gate_1957(n2033,n2032);
and gate_1958(n2034,n197,n2033);
not gate_1959(n2035,n2034);
and gate_1960(n2036,n2027,n2035);
not gate_1961(n2037,n2036);
and gate_1962(n2038,n84,n2037);
not gate_1963(n2039,n2038);
and gate_1964(n2040,n2025,n2039);
not gate_1965(n2041,n2040);
and gate_1966(n2042,n107,n2041);
and gate_1967(n2043,n104,n2042);
and gate_1968(n2044,n81,n2043);
not gate_1969(n2045,n2044);
and gate_1970(n2046,pi39,n126);
and gate_1971(n2047,n110,n2046);
and gate_1972(n2048,pi34,n2047);
not gate_1973(n2049,n2048);
and gate_1974(n2050,n2045,n2049);
not gate_1975(n2051,n2050);
and gate_1976(n2052,pi38,n2051);
not gate_1977(n2053,n2052);
and gate_1978(n2054,n90,n104);
and gate_1979(n2055,n84,n2054);
and gate_1980(n2056,n107,n2016);
and gate_1981(n2057,pi15,n2056);
and gate_1982(n2058,n2055,n2057);
and gate_1983(n2059,n81,n2058);
not gate_1984(n2060,n2059);
and gate_1985(n2061,n2053,n2060);
and gate_1986(n2062,n2015,n2061);
not gate_1987(n2063,n2062);
and gate_1988(n2064,n108,n2063);
not gate_1989(n2065,n2064);
and gate_1990(n2066,n182,n330);
not gate_1991(n2067,n2066);
and gate_1992(n2068,n110,n2067);
not gate_1993(n2069,n2068);
and gate_1994(n2070,n623,n2069);
not gate_1995(n2071,n2070);
and gate_1996(n2072,n758,n2071);
not gate_1997(n2073,n2072);
and gate_1998(n2074,n98,n324);
not gate_1999(n2075,n2074);
and gate_2000(n2076,n181,n1827);
not gate_2001(n2077,n2076);
and gate_2002(n2078,n2075,n2077);
not gate_2003(n2079,n2078);
and gate_2004(n2080,n110,n2079);
not gate_2005(n2081,n2080);
and gate_2006(n2082,n98,n373);
not gate_2007(n2083,n2082);
and gate_2008(n2084,n2081,n2083);
and gate_2009(n2085,n2073,n2084);
not gate_2010(n2086,n2085);
and gate_2011(n2087,n379,n2086);
and gate_2012(n2088,n197,n2087);
and gate_2013(n2089,n81,n2088);
not gate_2014(n2090,n2089);
and gate_2015(n2091,n2065,n2090);
not gate_2016(n2092,n2091);
and gate_2017(n2093,n109,n2092);
not gate_2018(n2094,n2093);
and gate_2019(n2095,n77,n114);
and gate_2020(n2096,pi04,n118);
and gate_2021(n2097,n2095,n2096);
not gate_2022(n2098,n2097);
and gate_2023(n2099,n137,n2098);
not gate_2024(n2100,n2099);
and gate_2025(n2101,pi38,n2100);
not gate_2026(n2102,n2101);
and gate_2027(n2103,n151,n2102);
not gate_2028(n2104,n2103);
and gate_2029(n2105,pi00,n2104);
not gate_2030(n2106,n2105);
and gate_2031(n2107,n118,n205);
not gate_2032(n2108,n2107);
and gate_2033(n2109,pi27,n108);
and gate_2034(n2110,pi10,n2109);
and gate_2035(n2111,n616,n2110);
not gate_2036(n2112,n2111);
and gate_2037(n2113,n2108,n2112);
not gate_2038(n2114,n2113);
and gate_2039(n2115,n113,n2114);
not gate_2040(n2116,n2115);
and gate_2041(n2117,n2106,n2116);
not gate_2042(n2118,n2117);
and gate_2043(n2119,n422,n2118);
not gate_2044(n2120,n2119);
and gate_2045(n2121,n2094,n2120);
not gate_2046(n2122,n2121);
and gate_2047(n2123,n105,n2122);
not gate_2048(n2124,n2123);
and gate_2049(n2125,n83,n2124);
not gate_2050(n2126,n2125);
and gate_2051(po17,pi33,n2126);
and gate_2052(n2128,n389,n671);
not gate_2053(n2129,n2128);
and gate_2054(n2130,n757,n1509);
and gate_2055(n2131,n486,n2130);
not gate_2056(n2132,n2131);
and gate_2057(n2133,n2129,n2132);
not gate_2058(n2134,n2133);
and gate_2059(n2135,n81,n2134);
not gate_2060(n2136,n2135);
and gate_2061(n2137,n157,n390);
not gate_2062(n2138,n2137);
and gate_2063(n2139,pi38,n2138);
not gate_2064(n2140,n2139);
and gate_2065(n2141,n2136,n2140);
not gate_2066(n2142,n2141);
and gate_2067(n2143,pi35,n2142);
not gate_2068(n2144,n2143);
and gate_2069(n2145,n125,n206);
and gate_2070(n2146,pi00,n2145);
not gate_2071(n2147,n2146);
and gate_2072(n2148,pi11,pi39);
not gate_2073(n2149,n2148);
and gate_2074(n2150,n111,n2149);
not gate_2075(n2151,n2150);
and gate_2076(n2152,n390,n2151);
and gate_2077(n2153,n2147,n2152);
not gate_2078(n2154,n2153);
and gate_2079(n2155,n1403,n2154);
not gate_2080(n2156,n2155);
and gate_2081(n2157,n2144,n2156);
not gate_2082(n2158,n2157);
and gate_2083(n2159,pi40,n2158);
not gate_2084(n2160,n2159);
and gate_2085(n2161,n110,n1736);
not gate_2086(n2162,n2161);
and gate_2087(n2163,n497,n2162);
not gate_2088(n2164,n2163);
and gate_2089(n2165,n109,n2164);
not gate_2090(n2166,n2165);
and gate_2091(n2167,n1598,n2166);
not gate_2092(n2168,n2167);
and gate_2093(n2169,n486,n757);
not gate_2094(n2170,n2169);
and gate_2095(n2171,n2168,n2169);
and gate_2096(n2172,n81,n2171);
not gate_2097(n2173,n2172);
and gate_2098(n2174,n1406,n1954);
not gate_2099(n2175,n2174);
and gate_2100(n2176,n1510,n2175);
not gate_2101(n2177,n2176);
and gate_2102(n2178,n112,n2177);
not gate_2103(n2179,n2178);
and gate_2104(n2180,pi36,n1076);
not gate_2105(n2181,n2180);
and gate_2106(n2182,pi38,n2181);
and gate_2107(n2183,pi00,n2182);
not gate_2108(n2184,n2183);
and gate_2109(n2185,n109,n957);
not gate_2110(n2186,n2185);
and gate_2111(n2187,n2184,n2186);
and gate_2112(n2188,n2179,n2187);
not gate_2113(n2189,n2188);
and gate_2114(n2190,pi37,n2189);
not gate_2115(n2191,n2190);
and gate_2116(n2192,n561,n2191);
and gate_2117(n2193,n2173,n2192);
not gate_2118(n2194,n2193);
and gate_2119(n2195,pi35,n2194);
not gate_2120(n2196,n2195);
and gate_2121(n2197,n112,n411);
not gate_2122(n2198,n2197);
and gate_2123(n2199,pi37,n2198);
not gate_2124(n2200,n2199);
and gate_2125(n2201,n112,n412);
not gate_2126(n2202,n2201);
and gate_2127(n2203,n410,n2202);
not gate_2128(n2204,n2203);
and gate_2129(n2205,n2200,n2204);
not gate_2130(n2206,n2205);
and gate_2131(n2207,n1403,n2206);
not gate_2132(n2208,n2207);
and gate_2133(n2209,n2196,n2208);
and gate_2134(n2210,n2160,n2209);
not gate_2135(n2211,n2210);
and gate_2136(n2212,n105,n2211);
not gate_2137(n2213,n2212);
and gate_2138(n2214,n220,n633);
not gate_2139(n2215,n2214);
and gate_2140(n2216,n647,n2215);
not gate_2141(n2217,n2216);
and gate_2142(n2218,n196,n255);
and gate_2143(n2219,n112,n2218);
not gate_2144(n2220,n2219);
and gate_2145(n2221,pi11,pi12);
not gate_2146(n2222,n2221);
and gate_2147(n2223,pi09,n2221);
not gate_2148(n2224,n2223);
and gate_2149(n2225,n2220,n2224);
not gate_2150(n2226,n2225);
and gate_2151(n2227,pi15,n2226);
not gate_2152(n2228,n2227);
and gate_2153(n2229,n131,n2228);
not gate_2154(n2230,n2229);
and gate_2155(n2231,n113,n2230);
not gate_2156(n2232,n2231);
and gate_2157(n2233,pi09,n988);
not gate_2158(n2234,n2233);
and gate_2159(n2235,n2232,n2234);
not gate_2160(n2236,n2235);
and gate_2161(n2237,pi38,n2236);
not gate_2162(n2238,n2237);
and gate_2163(n2239,pi37,n401);
not gate_2164(n2240,n2239);
and gate_2165(n2241,n2218,n2240);
and gate_2166(n2242,pi15,n2241);
not gate_2167(n2243,n2242);
and gate_2168(n2244,n825,n2243);
not gate_2169(n2245,n2244);
and gate_2170(n2246,n111,n2245);
not gate_2171(n2247,n2246);
and gate_2172(n2248,n2238,n2247);
and gate_2173(n2249,n2217,n2248);
not gate_2174(n2250,n2249);
and gate_2175(n2251,n104,n2250);
and gate_2176(n2252,n81,n2251);
not gate_2177(n2253,n2252);
and gate_2178(n2254,n653,n1145);
not gate_2179(n2255,n2254);
and gate_2180(n2256,n105,n2255);
and gate_2181(n2257,n2253,n2256);
not gate_2182(n2258,n2257);
and gate_2183(n2259,n170,n2258);
not gate_2184(n2260,n2259);
and gate_2185(n2261,n2213,n2260);
not gate_2186(n2262,n2261);
and gate_2187(n2263,n107,n2262);
not gate_2188(n2264,n2263);
and gate_2189(n2265,n81,n1668);
not gate_2190(n2266,n2265);
and gate_2191(n2267,pi37,n2266);
not gate_2192(n2268,n2267);
and gate_2193(n2269,n1173,n2268);
not gate_2194(n2270,n2269);
and gate_2195(n2271,n148,n2270);
not gate_2196(n2272,n2271);
and gate_2197(n2273,pi39,n2272);
not gate_2198(n2274,n2273);
and gate_2199(n2275,n194,n2274);
and gate_2200(n2276,n223,n390);
not gate_2201(n2277,n2276);
and gate_2202(n2278,pi00,n2277);
not gate_2203(n2279,n2278);
and gate_2204(n2280,n135,n411);
not gate_2205(n2281,n2280);
and gate_2206(n2282,n584,n2281);
not gate_2207(n2283,n2282);
and gate_2208(n2284,n2279,n2283);
not gate_2209(n2285,n2284);
and gate_2210(n2286,n1075,n2285);
not gate_2211(n2287,n2286);
and gate_2212(n2288,n2275,n2287);
not gate_2213(n2289,n2288);
and gate_2214(n2290,n1783,n2289);
not gate_2215(n2291,n2290);
and gate_2216(n2292,n600,n2291);
not gate_2217(n2293,n2292);
and gate_2218(n2294,n108,n2293);
and gate_2219(n2295,n105,n2294);
not gate_2220(n2296,n2295);
and gate_2221(n2297,n2264,n2296);
not gate_2222(n2298,n2297);
and gate_2223(n2299,pi33,n2298);
and gate_2224(po18,n83,n2299);
and gate_2225(n2301,n422,n1936);
not gate_2226(n2302,n2301);
and gate_2227(n2303,n110,n401);
and gate_2228(n2304,pi04,n2303);
and gate_2229(n2305,pi00,n2304);
not gate_2230(n2306,n2305);
and gate_2231(n2307,n130,n1252);
not gate_2232(n2308,n2307);
and gate_2233(n2309,n2306,n2308);
not gate_2234(n2310,n2309);
and gate_2235(n2311,n1783,n2310);
and gate_2236(n2312,n586,n2311);
not gate_2237(n2313,n2312);
and gate_2238(n2314,n2302,n2313);
not gate_2239(n2315,n2314);
and gate_2240(n2316,n108,n2315);
not gate_2241(n2317,n2316);
and gate_2242(n2318,n109,n128);
not gate_2243(n2319,n2318);
and gate_2244(n2320,n82,n112);
not gate_2245(n2321,n2320);
and gate_2246(n2322,pi36,pi37);
and gate_2247(n2323,n2321,n2322);
not gate_2248(n2324,n2323);
and gate_2249(n2325,n2319,n2324);
not gate_2250(n2326,n2325);
and gate_2251(n2327,n1461,n2326);
and gate_2252(n2328,n107,n2327);
not gate_2253(n2329,n2328);
and gate_2254(n2330,n2317,n2329);
not gate_2255(n2331,n2330);
and gate_2256(n2332,n111,n2331);
not gate_2257(n2333,n2332);
and gate_2258(n2334,n156,n1759);
not gate_2259(n2335,n2334);
and gate_2260(n2336,n379,n557);
not gate_2261(n2337,n2336);
and gate_2262(n2338,n2335,n2337);
not gate_2263(n2339,n2338);
and gate_2264(n2340,pi06,n400);
not gate_2265(n2341,n2340);
and gate_2266(n2342,n2339,n2340);
not gate_2267(n2343,n2342);
and gate_2268(n2344,pi00,n123);
and gate_2269(n2345,n143,n2322);
and gate_2270(n2346,n2344,n2345);
not gate_2271(n2347,n2346);
and gate_2272(n2348,n327,n1891);
not gate_2273(n2349,n2348);
and gate_2274(n2350,n2347,n2349);
not gate_2275(n2351,n2350);
and gate_2276(n2352,n379,n2351);
not gate_2277(n2353,n2352);
and gate_2278(n2354,n2343,n2353);
not gate_2279(n2355,n2354);
and gate_2280(n2356,pi38,n2355);
not gate_2281(n2357,n2356);
and gate_2282(n2358,n2333,n2357);
not gate_2283(n2359,n2358);
and gate_2284(po19,n429,n2359);
and gate_2285(n2361,pi35,n2067);
not gate_2286(n2362,n2361);
and gate_2287(n2363,n108,n218);
not gate_2288(n2364,n2363);
and gate_2289(n2365,n323,n2363);
not gate_2290(n2366,n2365);
and gate_2291(n2367,n84,n113);
not gate_2292(n2368,n2367);
and gate_2293(n2369,n181,n2368);
not gate_2294(n2370,n2369);
and gate_2295(n2371,n2366,n2370);
and gate_2296(n2372,n2362,n2371);
not gate_2297(n2373,n2372);
and gate_2298(n2374,n110,n2373);
not gate_2299(n2375,n2374);
and gate_2300(n2376,n108,n780);
not gate_2301(n2377,n2376);
and gate_2302(n2378,pi40,n1364);
not gate_2303(n2379,n2378);
and gate_2304(n2380,n2377,n2379);
not gate_2305(n2381,n2380);
and gate_2306(n2382,n185,n2381);
not gate_2307(n2383,n2382);
and gate_2308(n2384,n2375,n2383);
not gate_2309(n2385,n2384);
and gate_2310(n2386,n107,n2385);
not gate_2311(n2387,n2386);
and gate_2312(n2388,n1493,n1646);
not gate_2313(n2389,n2388);
and gate_2314(n2390,n2387,n2389);
not gate_2315(n2391,n2390);
and gate_2316(n2392,n198,n2391);
not gate_2317(n2393,n2392);
and gate_2318(n2394,n184,n374);
not gate_2319(n2395,n2394);
and gate_2320(n2396,pi35,n2395);
not gate_2321(n2397,n2396);
and gate_2322(n2398,n169,n1873);
not gate_2323(n2399,n2398);
and gate_2324(n2400,n112,n2399);
not gate_2325(n2401,n2400);
and gate_2326(n2402,n110,n805);
not gate_2327(n2403,n2402);
and gate_2328(n2404,n76,n113);
not gate_2329(n2405,n2404);
and gate_2330(n2406,n2403,n2405);
not gate_2331(n2407,n2406);
and gate_2332(n2408,pi39,n2407);
not gate_2333(n2409,n2408);
and gate_2334(n2410,n1494,n2409);
not gate_2335(n2411,n2410);
and gate_2336(n2412,pi38,n2411);
not gate_2337(n2413,n2412);
and gate_2338(n2414,n130,n802);
not gate_2339(n2415,n2414);
and gate_2340(n2416,n111,n2415);
and gate_2341(n2417,n108,n2416);
not gate_2342(n2418,n2417);
and gate_2343(n2419,n2413,n2418);
and gate_2344(n2420,n2401,n2419);
and gate_2345(n2421,n2397,n2420);
not gate_2346(n2422,n2421);
and gate_2347(n2423,pi05,n2422);
not gate_2348(n2424,n2423);
and gate_2349(n2425,n1136,n1138);
and gate_2350(n2426,n802,n2425);
not gate_2351(n2427,n2426);
and gate_2352(n2428,pi31,n2427);
not gate_2353(n2429,n2428);
and gate_2354(n2430,n190,n263);
not gate_2355(n2431,n2430);
and gate_2356(n2432,n881,n2431);
not gate_2357(n2433,n2432);
and gate_2358(n2434,pi09,n2433);
not gate_2359(n2435,n2434);
and gate_2360(n2436,n277,n651);
not gate_2361(n2437,n2436);
and gate_2362(n2438,n2435,n2437);
not gate_2363(n2439,n2438);
and gate_2364(n2440,n2222,n2439);
not gate_2365(n2441,n2440);
and gate_2366(n2442,n88,n652);
not gate_2367(n2443,n2442);
and gate_2368(n2444,n2441,n2443);
and gate_2369(n2445,n2429,n2444);
not gate_2370(n2446,n2445);
and gate_2371(n2447,n108,n2446);
not gate_2372(n2448,n2447);
and gate_2373(n2449,n2424,n2448);
not gate_2374(n2450,n2449);
and gate_2375(n2451,n107,n2450);
not gate_2376(n2452,n2451);
and gate_2377(n2453,n111,n2240);
not gate_2378(n2454,n2453);
and gate_2379(n2455,n76,n401);
not gate_2380(n2456,n2455);
and gate_2381(n2457,n110,n2456);
not gate_2382(n2458,n2457);
and gate_2383(n2459,n2453,n2458);
and gate_2384(n2460,n108,n2459);
and gate_2385(n2461,pi05,n2460);
not gate_2386(n2462,n2461);
and gate_2387(n2463,n2452,n2462);
and gate_2388(n2464,n2393,n2463);
not gate_2389(n2465,n2464);
and gate_2390(n2466,n109,n2465);
not gate_2391(n2467,n2466);
and gate_2392(n2468,n110,n205);
and gate_2393(n2469,n399,n2468);
not gate_2394(n2470,n2469);
and gate_2395(n2471,n108,n128);
not gate_2396(n2472,n2471);
and gate_2397(n2473,n131,n2472);
not gate_2398(n2474,n2473);
and gate_2399(n2475,pi38,n2474);
and gate_2400(n2476,n1885,n2475);
not gate_2401(n2477,n2476);
and gate_2402(n2478,n2470,n2477);
not gate_2403(n2479,n2478);
and gate_2404(n2480,pi40,n2479);
not gate_2405(n2481,n2480);
and gate_2406(n2482,pi35,n535);
and gate_2407(n2483,n1885,n2482);
not gate_2408(n2484,n2483);
and gate_2409(n2485,n2481,n2484);
not gate_2410(n2486,n2485);
and gate_2411(n2487,n422,n2486);
not gate_2412(n2488,n2487);
and gate_2413(n2489,n2467,n2488);
not gate_2414(n2490,n2489);
and gate_2415(po20,n429,n2490);
and gate_2416(n2492,n81,pi38);
not gate_2417(n2493,n2492);
and gate_2418(n2494,n330,n2493);
not gate_2419(n2495,n2494);
and gate_2420(n2496,n76,n2495);
not gate_2421(n2497,n2496);
and gate_2422(n2498,n1173,n2320);
not gate_2423(n2499,n2498);
and gate_2424(n2500,n2497,n2499);
not gate_2425(n2501,n2500);
and gate_2426(n2502,pi37,n2501);
not gate_2427(n2503,n2502);
and gate_2428(n2504,n82,n449);
not gate_2429(n2505,n2504);
and gate_2430(n2506,n2503,n2505);
not gate_2431(n2507,n2506);
and gate_2432(n2508,pi35,n2507);
not gate_2433(n2509,n2508);
and gate_2434(n2510,n1303,n2474);
and gate_2435(n2511,n81,n2510);
and gate_2436(n2512,n76,n2511);
not gate_2437(n2513,n2512);
and gate_2438(n2514,n105,n2513);
and gate_2439(n2515,n2509,n2514);
not gate_2440(n2516,n2515);
and gate_2441(n2517,pi36,n2516);
not gate_2442(n2518,n2517);
and gate_2443(n2519,n76,n1046);
and gate_2444(n2520,n161,n2519);
not gate_2445(n2521,n2520);
and gate_2446(n2522,n105,n2521);
not gate_2447(n2523,n2522);
and gate_2448(n2524,pi35,n2523);
not gate_2449(n2525,n2524);
and gate_2450(n2526,n2518,n2525);
not gate_2451(n2527,n2526);
and gate_2452(n2528,n107,n2527);
not gate_2453(n2529,n2528);
and gate_2454(n2530,n110,n1753);
and gate_2455(n2531,n81,n2530);
and gate_2456(n2532,n76,n2531);
not gate_2457(n2533,n2532);
and gate_2458(n2534,n82,pi37);
and gate_2459(n2535,n703,n2534);
not gate_2460(n2536,n2535);
and gate_2461(n2537,n105,n2536);
and gate_2462(n2538,n2533,n2537);
not gate_2463(n2539,n2538);
and gate_2464(n2540,n1783,n2539);
not gate_2465(n2541,n2540);
and gate_2466(n2542,pi32,n599);
not gate_2467(n2543,n2542);
and gate_2468(n2544,n2541,n2543);
not gate_2469(n2545,n2544);
and gate_2470(n2546,n108,n2545);
not gate_2471(n2547,n2546);
and gate_2472(n2548,n2529,n2547);
not gate_2473(n2549,n2548);
and gate_2474(n2550,n83,n2549);
not gate_2475(n2551,n2550);
and gate_2476(n2552,pi33,n2551);
not gate_2477(po21,n2552);
and gate_2478(n2554,n263,n2221);
and gate_2479(n2555,n510,n2554);
and gate_2480(n2556,n2425,n2555);
and gate_2481(n2557,n432,n2556);
not gate_2482(n2558,n2557);
and gate_2483(n2559,pi05,n2558);
not gate_2484(n2560,n2559);
and gate_2485(n2561,n527,n2454);
not gate_2486(n2562,n2561);
and gate_2487(n2563,n2218,n2562);
not gate_2488(n2564,n2563);
and gate_2489(n2565,n779,n2223);
not gate_2490(n2566,n2565);
and gate_2491(n2567,n2564,n2566);
not gate_2492(n2568,n2567);
and gate_2493(n2569,pi15,n2568);
not gate_2494(n2570,n2569);
and gate_2495(n2571,n327,n1578);
not gate_2496(n2572,n2571);
and gate_2497(n2573,n2570,n2572);
not gate_2498(n2574,n2573);
and gate_2499(n2575,n104,n2574);
not gate_2500(n2576,n2575);
and gate_2501(n2577,n105,n2576);
and gate_2502(n2578,n2560,n2577);
not gate_2503(n2579,n2578);
and gate_2504(n2580,n108,n2579);
not gate_2505(n2581,n2580);
and gate_2506(n2582,n1598,n2397);
not gate_2507(n2583,n2582);
and gate_2508(n2584,n105,n2583);
and gate_2509(n2585,pi05,n2584);
not gate_2510(n2586,n2585);
and gate_2511(n2587,n2581,n2586);
not gate_2512(n2588,n2587);
and gate_2513(n2589,n109,n2588);
not gate_2514(n2590,n2589);
and gate_2515(n2591,n109,n160);
not gate_2516(n2592,n2591);
and gate_2517(n2593,pi35,n2591);
not gate_2518(n2594,n2593);
and gate_2519(n2595,n2364,n2594);
and gate_2520(n2596,pi37,n2595);
not gate_2521(n2597,n2596);
and gate_2522(n2598,n402,n1403);
not gate_2523(n2599,n2598);
and gate_2524(n2600,n2597,n2599);
not gate_2525(n2601,n2600);
and gate_2526(n2602,pi38,n2601);
and gate_2527(n2603,n105,n2602);
and gate_2528(n2604,n1885,n2603);
not gate_2529(n2605,n2604);
and gate_2530(n2606,n2590,n2605);
not gate_2531(n2607,n2606);
and gate_2532(n2608,n107,n2607);
not gate_2533(n2609,n2608);
and gate_2534(n2610,n170,n2459);
and gate_2535(n2611,n105,n2610);
and gate_2536(n2612,pi05,n2611);
not gate_2537(n2613,n2612);
and gate_2538(n2614,n2609,n2613);
not gate_2539(n2615,n2614);
and gate_2540(n2616,pi33,n2615);
and gate_2541(po22,n83,n2616);
and gate_2542(n2618,n107,n535);
not gate_2543(n2619,n2618);
and gate_2544(n2620,n172,n2619);
not gate_2545(n2621,n2620);
and gate_2546(n2622,n76,n2621);
not gate_2547(n2623,n2622);
and gate_2548(n2624,pi36,n111);
not gate_2549(n2625,n2624);
and gate_2550(n2626,n107,n108);
and gate_2551(n2627,n2625,n2626);
not gate_2552(n2628,n2627);
and gate_2553(n2629,n2623,n2628);
not gate_2554(n2630,n2629);
and gate_2555(n2631,pi05,n2630);
not gate_2556(n2632,n2631);
and gate_2557(n2633,n1888,n1894);
not gate_2558(n2634,n2633);
and gate_2559(n2635,n80,n2634);
not gate_2560(n2636,n2635);
and gate_2561(n2637,n111,n1686);
not gate_2562(n2638,n2637);
and gate_2563(n2639,n1888,n2638);
not gate_2564(n2640,n2639);
and gate_2565(n2641,n114,n2640);
not gate_2566(n2642,n2641);
and gate_2567(n2643,n2636,n2642);
not gate_2568(n2644,n2643);
and gate_2569(n2645,n77,n2644);
not gate_2570(n2646,n2645);
and gate_2571(n2647,n108,n1435);
not gate_2572(n2648,n2647);
and gate_2573(n2649,pi36,n1407);
not gate_2574(n2650,n2649);
and gate_2575(n2651,n118,n2650);
not gate_2576(n2652,n2651);
and gate_2577(n2653,n2648,n2652);
not gate_2578(n2654,n2653);
and gate_2579(n2655,n107,n2654);
not gate_2580(n2656,n2655);
and gate_2581(n2657,n2646,n2656);
not gate_2582(n2658,n2657);
and gate_2583(n2659,pi00,n2658);
not gate_2584(n2660,n2659);
and gate_2585(n2661,n109,pi39);
not gate_2586(n2662,n2661);
and gate_2587(n2663,n113,n2662);
not gate_2588(n2664,n2663);
and gate_2589(n2665,n111,n2664);
and gate_2590(n2666,n107,n2665);
not gate_2591(n2667,n2666);
and gate_2592(n2668,n109,n447);
not gate_2593(n2669,n2668);
and gate_2594(n2670,n2667,n2669);
not gate_2595(n2671,n2670);
and gate_2596(n2672,n198,n2671);
not gate_2597(n2673,n2672);
and gate_2598(n2674,n1174,n2662);
not gate_2599(n2675,n2674);
and gate_2600(n2676,n90,n2675);
not gate_2601(n2677,n2676);
and gate_2602(n2678,n109,n181);
not gate_2603(n2679,n2678);
and gate_2604(n2680,n2677,n2679);
not gate_2605(n2681,n2680);
and gate_2606(n2682,n84,n2681);
not gate_2607(n2683,n2682);
and gate_2608(n2684,pi38,n1203);
not gate_2609(n2685,n2684);
and gate_2610(n2686,n989,n1174);
and gate_2611(n2687,n2685,n2686);
not gate_2612(n2688,n2687);
and gate_2613(n2689,pi36,n2688);
not gate_2614(n2690,n2689);
and gate_2615(n2691,pi31,n109);
not gate_2616(n2692,n2691);
and gate_2617(n2693,n2690,n2692);
and gate_2618(n2694,n2683,n2693);
not gate_2619(n2695,n2694);
and gate_2620(n2696,n107,n2695);
not gate_2621(n2697,n2696);
and gate_2622(n2698,pi34,n1509);
not gate_2623(n2699,n2698);
and gate_2624(n2700,n185,n557);
not gate_2625(n2701,n2700);
and gate_2626(n2702,n2699,n2701);
not gate_2627(n2703,n2702);
and gate_2628(n2704,n113,n2703);
not gate_2629(n2705,n2704);
and gate_2630(n2706,n107,n113);
not gate_2631(n2707,n2706);
and gate_2632(n2708,n989,n2707);
not gate_2633(n2709,n2708);
and gate_2634(n2710,pi39,n2222);
not gate_2635(n2711,n2710);
and gate_2636(n2712,n255,n2711);
not gate_2637(n2713,n2712);
and gate_2638(n2714,n110,n2713);
not gate_2639(n2715,n2714);
and gate_2640(n2716,n2709,n2715);
not gate_2641(n2717,n2716);
and gate_2642(n2718,pi38,n2717);
not gate_2643(n2719,n2718);
and gate_2644(n2720,n113,n125);
not gate_2645(n2721,n2720);
and gate_2646(n2722,pi37,n2721);
not gate_2647(n2723,n2722);
and gate_2648(n2724,n1975,n2723);
not gate_2649(n2725,n2724);
and gate_2650(n2726,n111,n2725);
and gate_2651(n2727,pi34,n2726);
not gate_2652(n2728,n2727);
and gate_2653(n2729,n2719,n2728);
not gate_2654(n2730,n2729);
and gate_2655(n2731,n109,n2730);
not gate_2656(n2732,n2731);
and gate_2657(n2733,n2705,n2732);
and gate_2658(n2734,n2697,n2733);
and gate_2659(n2735,n2673,n2734);
not gate_2660(n2736,n2735);
and gate_2661(n2737,n108,n2736);
not gate_2662(n2738,n2737);
and gate_2663(n2739,pi38,n1085);
not gate_2664(n2740,n2739);
and gate_2665(n2741,n111,n2662);
not gate_2666(n2742,n2741);
and gate_2667(n2743,n218,n2742);
and gate_2668(n2744,n2740,n2743);
not gate_2669(n2745,n2744);
and gate_2670(n2746,n110,n2745);
not gate_2671(n2747,n2746);
and gate_2672(n2748,n223,n2592);
not gate_2673(n2749,n2748);
and gate_2674(n2750,pi37,n2749);
not gate_2675(n2751,n2750);
and gate_2676(n2752,n2747,n2751);
not gate_2677(n2753,n2752);
and gate_2678(n2754,pi35,n2753);
not gate_2679(n2755,n2754);
and gate_2680(n2756,n156,n1753);
not gate_2681(n2757,n2756);
and gate_2682(n2758,n2755,n2757);
not gate_2683(n2759,n2758);
and gate_2684(n2760,n107,n2759);
not gate_2685(n2761,n2760);
and gate_2686(n2762,n2738,n2761);
and gate_2687(n2763,n2660,n2762);
and gate_2688(n2764,n2632,n2763);
not gate_2689(n2765,n2764);
and gate_2690(n2766,n105,n2765);
not gate_2691(n2767,n2766);
and gate_2692(n2768,n83,n2767);
not gate_2693(n2769,n2768);
and gate_2694(po23,pi33,n2769);
and gate_2695(n2771,n126,n133);
and gate_2696(n2772,pi36,n2771);
and gate_2697(n2773,pi00,n2772);
not gate_2698(n2774,n2773);
and gate_2699(n2775,n109,n2023);
and gate_2700(n2776,n104,n2775);
and gate_2701(n2777,n81,n2776);
not gate_2702(n2778,n2777);
and gate_2703(n2779,n2774,n2778);
not gate_2704(n2780,n2779);
and gate_2705(n2781,pi40,n2780);
not gate_2706(n2782,n2781);
and gate_2707(n2783,n104,n109);
and gate_2708(n2784,n2038,n2783);
and gate_2709(n2785,n81,n2784);
not gate_2710(n2786,n2785);
and gate_2711(n2787,pi36,n824);
and gate_2712(n2788,n412,n2787);
not gate_2713(n2789,n2788);
and gate_2714(n2790,n2786,n2789);
and gate_2715(n2791,n2782,n2790);
not gate_2716(n2792,n2791);
and gate_2717(n2793,pi38,n2792);
not gate_2718(n2794,n2793);
and gate_2719(n2795,n111,n1276);
not gate_2720(n2796,n2795);
and gate_2721(n2797,n128,n254);
not gate_2722(n2798,n2797);
and gate_2723(n2799,n2796,n2798);
not gate_2724(n2800,n2799);
and gate_2725(n2801,n197,n2800);
not gate_2726(n2802,n2801);
and gate_2727(n2803,n496,n1995);
not gate_2728(n2804,n2803);
and gate_2729(n2805,n2802,n2804);
not gate_2730(n2806,n2805);
and gate_2731(n2807,n2783,n2806);
and gate_2732(n2808,n81,n2807);
not gate_2733(n2809,n2808);
and gate_2734(n2810,n2794,n2809);
not gate_2735(n2811,n2810);
and gate_2736(n2812,n108,n2811);
not gate_2737(n2813,n2812);
and gate_2738(n2814,n1006,n1407);
not gate_2739(n2815,n2814);
and gate_2740(n2816,n77,n2815);
not gate_2741(n2817,n2816);
and gate_2742(n2818,n78,n143);
not gate_2743(n2819,n2818);
and gate_2744(n2820,n1406,n2819);
not gate_2745(n2821,n2820);
and gate_2746(n2822,n2817,n2821);
not gate_2747(n2823,n2822);
and gate_2748(n2824,pi00,n2823);
not gate_2749(n2825,n2824);
and gate_2750(n2826,n223,n2825);
not gate_2751(n2827,n2826);
and gate_2752(n2828,pi36,n2827);
not gate_2753(n2829,n2828);
and gate_2754(n2830,n95,n362);
not gate_2755(n2831,n2830);
and gate_2756(n2832,pi22,n2831);
not gate_2757(n2833,n2832);
and gate_2758(n2834,n1697,n2833);
and gate_2759(n2835,n111,n2834);
and gate_2760(n2836,pi15,n2835);
and gate_2761(n2837,n81,n2836);
not gate_2762(n2838,n2837);
and gate_2763(n2839,n411,n2838);
not gate_2764(n2840,n2839);
and gate_2765(n2841,n112,n2840);
and gate_2766(n2842,n109,n2841);
not gate_2767(n2843,n2842);
and gate_2768(n2844,n2829,n2843);
not gate_2769(n2845,n2844);
and gate_2770(n2846,pi37,n2845);
not gate_2771(n2847,n2846);
and gate_2772(n2848,n96,n2067);
not gate_2773(n2849,n2848);
and gate_2774(n2850,n95,n113);
not gate_2775(n2851,n2850);
and gate_2776(n2852,pi24,n2851);
not gate_2777(n2853,n2852);
and gate_2778(n2854,n324,n2853);
not gate_2779(n2855,n2854);
and gate_2780(n2856,n946,n1828);
not gate_2781(n2857,n2856);
and gate_2782(n2858,n181,n2857);
not gate_2783(n2859,n2858);
and gate_2784(n2860,n2855,n2859);
and gate_2785(n2861,n2849,n2860);
not gate_2786(n2862,n2861);
and gate_2787(n2863,n110,n2862);
not gate_2788(n2864,n2863);
and gate_2789(n2865,n2083,n2864);
not gate_2790(n2866,n2865);
and gate_2791(n2867,n109,n2866);
and gate_2792(n2868,n197,n2867);
and gate_2793(n2869,n81,n2868);
not gate_2794(n2870,n2869);
and gate_2795(n2871,n2847,n2870);
not gate_2796(n2872,n2871);
and gate_2797(n2873,pi35,n2872);
not gate_2798(n2874,n2873);
and gate_2799(n2875,n2813,n2874);
not gate_2800(n2876,n2875);
and gate_2801(n2877,n107,n2876);
not gate_2802(n2878,n2877);
and gate_2803(n2879,n111,n1992);
not gate_2804(n2880,n2879);
and gate_2805(n2881,n447,n2046);
not gate_2806(n2882,n2881);
and gate_2807(n2883,n2880,n2882);
not gate_2808(n2884,n2883);
and gate_2809(n2885,n109,n2884);
not gate_2810(n2886,n2885);
and gate_2811(n2887,n600,n2886);
not gate_2812(n2888,n2887);
and gate_2813(n2889,n1759,n2888);
not gate_2814(n2890,n2889);
and gate_2815(n2891,n2878,n2890);
not gate_2816(n2892,n2891);
and gate_2817(po24,n429,n2892);
and gate_2818(n2894,n2095,n2305);
not gate_2819(n2895,n2894);
and gate_2820(n2896,n1046,n1249);
not gate_2821(n2897,n2896);
and gate_2822(n2898,n2895,n2897);
not gate_2823(n2899,n2898);
and gate_2824(n2900,pi34,n2899);
not gate_2825(n2901,n2900);
and gate_2826(n2902,n2011,n2901);
not gate_2827(n2903,n2902);
and gate_2828(n2904,n108,n2903);
not gate_2829(n2905,n2904);
and gate_2830(n2906,pi37,n2833);
not gate_2831(n2907,n2906);
and gate_2832(n2908,pi24,n2907);
not gate_2833(n2909,n2908);
and gate_2834(n2910,pi40,n2909);
not gate_2835(n2911,n2910);
and gate_2836(n2912,n113,n758);
not gate_2837(n2913,n2912);
and gate_2838(n2914,pi24,n2913);
not gate_2839(n2915,n2914);
and gate_2840(n2916,n110,n2915);
not gate_2841(n2917,n2916);
and gate_2842(n2918,n2911,n2917);
not gate_2843(n2919,n2918);
and gate_2844(n2920,n112,n2919);
and gate_2845(n2921,n379,n2920);
and gate_2846(n2922,n197,n2921);
and gate_2847(n2923,n81,n2922);
not gate_2848(n2924,n2923);
and gate_2849(n2925,n2905,n2924);
not gate_2850(n2926,n2925);
and gate_2851(n2927,n111,n2926);
not gate_2852(n2928,n2927);
and gate_2853(n2929,n84,n2026);
not gate_2854(n2930,n2929);
and gate_2855(n2931,n217,n236);
not gate_2856(n2932,n2931);
and gate_2857(n2933,n2930,n2932);
not gate_2858(n2934,n2933);
and gate_2859(n2935,n1872,n2934);
and gate_2860(n2936,n104,n2935);
not gate_2861(n2937,n2936);
and gate_2862(n2938,n262,n275);
not gate_2863(n2939,n2938);
and gate_2864(n2940,n432,n2939);
not gate_2865(n2941,n2940);
and gate_2866(n2942,n108,n2941);
and gate_2867(n2943,n104,n2942);
not gate_2868(n2944,n2943);
and gate_2869(n2945,n95,n691);
not gate_2870(n2946,n2945);
and gate_2871(n2947,pi24,n1828);
and gate_2872(n2948,pi22,n2947);
and gate_2873(n2949,n2946,n2948);
not gate_2874(n2950,n2949);
and gate_2875(n2951,n547,n2950);
not gate_2876(n2952,n2951);
and gate_2877(n2953,n2944,n2952);
not gate_2878(n2954,n2953);
and gate_2879(n2955,pi39,n2954);
not gate_2880(n2956,n2955);
and gate_2881(n2957,n108,n779);
and gate_2882(n2958,n2055,n2957);
not gate_2883(n2959,n2958);
and gate_2884(n2960,n2956,n2959);
not gate_2885(n2961,n2960);
and gate_2886(n2962,pi38,n2961);
not gate_2887(n2963,n2962);
and gate_2888(n2964,n2055,n2471);
not gate_2889(n2965,n2964);
and gate_2890(n2966,n2963,n2965);
not gate_2891(n2967,n2966);
and gate_2892(n2968,n197,n2967);
not gate_2893(n2969,n2968);
and gate_2894(n2970,n2937,n2969);
not gate_2895(n2971,n2970);
and gate_2896(n2972,n107,n2971);
and gate_2897(n2973,n81,n2972);
not gate_2898(n2974,n2973);
and gate_2899(n2975,n2928,n2974);
not gate_2900(n2976,n2975);
and gate_2901(n2977,n109,n2976);
not gate_2902(n2978,n2977);
and gate_2903(n2979,n572,n2110);
not gate_2904(n2980,n2979);
and gate_2905(n2981,n79,n1004);
and gate_2906(n2982,pi02,n2981);
and gate_2907(n2983,n789,n2982);
not gate_2908(n2984,n2983);
and gate_2909(n2985,n223,n2984);
not gate_2910(n2986,n2985);
and gate_2911(n2987,n118,n2986);
not gate_2912(n2988,n2987);
and gate_2913(n2989,n2980,n2988);
not gate_2914(n2990,n2989);
and gate_2915(n2991,n107,n2990);
not gate_2916(n2992,n2991);
and gate_2917(n2993,pi34,n1621);
and gate_2918(n2994,n329,n2993);
not gate_2919(n2995,n2994);
and gate_2920(n2996,n2992,n2995);
not gate_2921(n2997,n2996);
and gate_2922(n2998,pi36,n2997);
not gate_2923(n2999,n2998);
and gate_2924(n3000,n2978,n2999);
not gate_2925(n3001,n3000);
and gate_2926(po25,n429,n3001);
and gate_2927(n3003,n134,n422);
and gate_2928(n3004,pi00,n3003);
not gate_2929(n3005,n3004);
and gate_2930(n3006,n128,n1783);
not gate_2931(n3007,n3006);
and gate_2932(n3008,n3005,n3007);
not gate_2933(n3009,n3008);
and gate_2934(n3010,pi38,n3009);
not gate_2935(n3011,n3010);
and gate_2936(n3012,n187,n1783);
not gate_2937(n3013,n3012);
and gate_2938(n3014,n3011,n3013);
not gate_2939(n3015,n3014);
and gate_2940(n3016,n126,n3015);
not gate_2941(n3017,n3016);
and gate_2942(n3018,n602,n3017);
not gate_2943(n3019,n3018);
and gate_2944(n3020,n108,n3019);
not gate_2945(n3021,n3020);
and gate_2946(n3022,n107,n1454);
and gate_2947(n3023,n146,n1936);
and gate_2948(n3024,n3022,n3023);
and gate_2949(n3025,pi00,n3024);
not gate_2950(n3026,n3025);
and gate_2951(n3027,n3021,n3026);
not gate_2952(n3028,n3027);
and gate_2953(po26,n429,n3028);
and gate_2954(n3030,n1872,n2026);
and gate_2955(n3031,n107,n3030);
and gate_2956(n3032,n104,n3031);
and gate_2957(n3033,n84,n3032);
not gate_2958(n3034,n3033);
and gate_2959(n3035,n111,n2920);
not gate_2960(n3036,n3035);
and gate_2961(n3037,n183,n2950);
not gate_2962(n3038,n3037);
and gate_2963(n3039,n3036,n3038);
not gate_2964(n3040,n3039);
and gate_2965(n3041,pi35,n3040);
not gate_2966(n3042,n3041);
and gate_2967(n3043,n91,n651);
not gate_2968(n3044,n3043);
and gate_2969(n3045,n110,n2198);
not gate_2970(n3046,n3045);
and gate_2971(n3047,n182,n293);
and gate_2972(n3048,n3046,n3047);
not gate_2973(n3049,n3048);
and gate_2974(n3050,n84,n3049);
not gate_2975(n3051,n3050);
and gate_2976(n3052,n3044,n3051);
not gate_2977(n3053,n3052);
and gate_2978(n3054,n90,n3053);
not gate_2979(n3055,n3054);
and gate_2980(n3056,n182,n188);
not gate_2981(n3057,n3056);
and gate_2982(n3058,n91,n3057);
and gate_2983(n3059,n84,n3058);
not gate_2984(n3060,n3059);
and gate_2985(n3061,n3055,n3060);
not gate_2986(n3062,n3061);
and gate_2987(n3063,n108,n3062);
and gate_2988(n3064,n104,n3063);
not gate_2989(n3065,n3064);
and gate_2990(n3066,n3042,n3065);
not gate_2991(n3067,n3066);
and gate_2992(n3068,n107,n3067);
not gate_2993(n3069,n3068);
and gate_2994(n3070,n614,n1247);
and gate_2995(n3071,n1759,n3070);
not gate_2996(n3072,n3071);
and gate_2997(n3073,n3069,n3072);
not gate_2998(n3074,n3073);
and gate_2999(n3075,n197,n3074);
not gate_3000(n3076,n3075);
and gate_3001(n3077,n3034,n3076);
not gate_3002(n3078,n3077);
and gate_3003(n3079,n109,n3078);
and gate_3004(n3080,n81,n3079);
not gate_3005(n3081,n3080);
and gate_3006(n3082,n632,n3022);
not gate_3007(n3083,n3082);
and gate_3008(n3084,n3081,n3083);
not gate_3009(n3085,n3084);
and gate_3010(po27,n429,n3085);
and gate_3011(n3087,n412,n2626);
and gate_3012(n3088,n526,n557);
and gate_3013(n3089,n3087,n3088);
not gate_3014(n3090,n3089);
and gate_3015(n3091,n1686,n2530);
not gate_3016(n3092,n3091);
and gate_3017(n3093,n1890,n3092);
not gate_3018(n3094,n3093);
and gate_3019(n3095,n783,n3094);
and gate_3020(n3096,n789,n3095);
not gate_3021(n3097,n3096);
and gate_3022(n3098,n3090,n3097);
not gate_3023(n3099,n3098);
and gate_3024(po28,n429,n3099);
and gate_3025(n3101,n324,n547);
and gate_3026(n3102,n692,n3101);
and gate_3027(n3103,n95,n3102);
and gate_3028(n3104,pi15,n3103);
not gate_3029(n3105,n3104);
and gate_3030(n3106,n236,n614);
and gate_3031(n3107,n108,n3106);
and gate_3032(n3108,n104,n3107);
not gate_3033(n3109,n3108);
and gate_3034(n3110,n3105,n3109);
not gate_3035(n3111,n3110);
and gate_3036(n3112,n113,n3111);
not gate_3037(n3113,n3112);
and gate_3038(n3114,n1872,n2931);
and gate_3039(n3115,n104,n3114);
not gate_3040(n3116,n3115);
and gate_3041(n3117,n3113,n3116);
not gate_3042(n3118,n3117);
and gate_3043(n3119,n107,n3118);
not gate_3044(n3120,n3119);
and gate_3045(n3121,n111,n1698);
not gate_3046(n3122,n3121);
and gate_3047(n3123,n1493,n3121);
and gate_3048(n3124,pi34,n3123);
and gate_3049(n3125,n341,n3124);
and gate_3050(n3126,pi15,n3125);
not gate_3051(n3127,n3126);
and gate_3052(n3128,n3120,n3127);
not gate_3053(n3129,n3128);
and gate_3054(n3130,n109,n3129);
and gate_3055(n3131,n81,n3130);
not gate_3056(n3132,n3131);
and gate_3057(n3133,n3083,n3132);
not gate_3058(n3134,n3133);
and gate_3059(po29,n429,n3134);
and gate_3060(n3136,pi37,n677);
and gate_3061(n3137,n97,n3136);
and gate_3062(n3138,pi40,n3137);
not gate_3063(n3139,n3138);
and gate_3064(n3140,n780,n3139);
not gate_3065(n3141,n3140);
and gate_3066(n3142,n95,n3141);
not gate_3067(n3143,n3142);
and gate_3068(n3144,n780,n1106);
not gate_3069(n3145,n3144);
and gate_3070(n3146,n96,n3145);
not gate_3071(n3147,n3146);
and gate_3072(n3148,n3143,n3147);
not gate_3073(n3149,n3148);
and gate_3074(n3150,n185,n3149);
not gate_3075(n3151,n3150);
and gate_3076(n3152,n113,n1030);
not gate_3077(n3153,n3152);
and gate_3078(n3154,pi22,n3153);
not gate_3079(n3155,n3154);
and gate_3080(n3156,n183,n3155);
not gate_3081(n3157,n3156);
and gate_3082(n3158,n3151,n3157);
not gate_3083(n3159,n3158);
and gate_3084(n3160,n379,n3159);
and gate_3085(n3161,pi24,n3160);
not gate_3086(n3162,n3161);
and gate_3087(n3163,n3072,n3162);
not gate_3088(n3164,n3163);
and gate_3089(n3165,n109,n3164);
and gate_3090(n3166,n197,n3165);
and gate_3091(n3167,n81,n3166);
not gate_3092(n3168,n3167);
and gate_3093(n3169,n3090,n3168);
not gate_3094(n3170,n3169);
and gate_3095(po30,n429,n3170);
and gate_3096(n3172,n98,n148);
not gate_3097(n3173,n3172);
and gate_3098(n3174,n341,n3137);
and gate_3099(n3175,pi40,n3174);
not gate_3100(n3176,n3175);
and gate_3101(n3177,n3173,n3176);
not gate_3102(n3178,n3177);
and gate_3103(n3179,n185,n3178);
not gate_3104(n3180,n3179);
and gate_3105(n3181,n757,n1827);
not gate_3106(n3182,n3181);
and gate_3107(n3183,pi24,n3182);
not gate_3108(n3184,n3183);
and gate_3109(n3185,n183,n3184);
not gate_3110(n3186,n3185);
and gate_3111(n3187,n3180,n3186);
not gate_3112(n3188,n3187);
and gate_3113(n3189,n109,n3188);
and gate_3114(n3190,n197,n3189);
and gate_3115(n3191,n81,n3190);
not gate_3116(n3192,n3191);
and gate_3117(n3193,n789,n2322);
and gate_3118(n3194,n1005,n3193);
not gate_3119(n3195,n3194);
and gate_3120(n3196,n3192,n3195);
not gate_3121(n3197,n3196);
and gate_3122(n3198,pi35,n3197);
not gate_3123(n3199,n3198);
and gate_3124(n3200,n412,n1403);
and gate_3125(n3201,n572,n3200);
not gate_3126(n3202,n3201);
and gate_3127(n3203,n3199,n3202);
not gate_3128(n3204,n3203);
and gate_3129(n3205,n107,n3204);
not gate_3130(n3206,n3205);
and gate_3131(n3207,n783,n3091);
and gate_3132(n3208,n789,n3207);
not gate_3133(n3209,n3208);
and gate_3134(n3210,n3206,n3209);
not gate_3135(n3211,n3210);
and gate_3136(po31,n429,n3211);
and gate_3137(n3213,n379,n429);
and gate_3138(n3214,n156,n3213);
and gate_3139(po32,n526,n3214);
and gate_3140(n3216,pi04,n110);
and gate_3141(n3217,pi00,n3216);
not gate_3142(n3218,n3217);
and gate_3143(n3219,n2308,n3218);
not gate_3144(n3220,n3219);
and gate_3145(n3221,n586,n3220);
not gate_3146(n3222,n3221);
and gate_3147(n3223,pi37,n1673);
not gate_3148(n3224,n3223);
and gate_3149(n3225,n400,n3224);
not gate_3150(n3226,n3225);
and gate_3151(n3227,n3222,n3226);
not gate_3152(n3228,n3227);
and gate_3153(n3229,pi34,n3228);
not gate_3154(n3230,n3229);
and gate_3155(n3231,n129,n290);
not gate_3156(n3232,n3231);
and gate_3157(n3233,n198,n3232);
not gate_3158(n3234,n3233);
and gate_3159(n3235,n443,n1146);
not gate_3160(n3236,n3235);
and gate_3161(n3237,n112,n3235);
not gate_3162(n3238,n3237);
and gate_3163(n3239,n159,n897);
not gate_3164(n3240,n3239);
and gate_3165(n3241,n3238,n3240);
not gate_3166(n3242,n3241);
and gate_3167(n3243,pi37,n3242);
not gate_3168(n3244,n3243);
and gate_3169(n3245,n3234,n3244);
not gate_3170(n3246,n3245);
and gate_3171(n3247,n107,n3246);
and gate_3172(n3248,n104,n3247);
and gate_3173(n3249,n81,n3248);
not gate_3174(n3250,n3249);
and gate_3175(n3251,n3230,n3250);
not gate_3176(n3252,n3251);
and gate_3177(n3253,n111,n3252);
not gate_3178(n3254,n3253);
and gate_3179(n3255,n107,n400);
not gate_3180(n3256,n3255);
and gate_3181(n3257,n527,n3256);
not gate_3182(n3258,n3257);
and gate_3183(n3259,n198,n3258);
not gate_3184(n3260,n3259);
and gate_3185(n3261,n703,n1146);
and gate_3186(n3262,n107,n3261);
and gate_3187(n3263,n277,n3262);
not gate_3188(n3264,n3263);
and gate_3189(n3265,n3260,n3264);
not gate_3190(n3266,n3265);
and gate_3191(n3267,n110,n3266);
not gate_3192(n3268,n3267);
and gate_3193(n3269,n88,pi40);
not gate_3194(n3270,n3269);
and gate_3195(n3271,n2221,n3270);
not gate_3196(n3272,n3271);
and gate_3197(n3273,n263,n3272);
not gate_3198(n3274,n3273);
and gate_3199(n3275,n110,n3274);
not gate_3200(n3276,n3275);
and gate_3201(n3277,n1297,n3276);
and gate_3202(n3278,pi09,n3277);
not gate_3203(n3279,n3278);
and gate_3204(n3280,n217,n897);
not gate_3205(n3281,n3280);
and gate_3206(n3282,n3279,n3281);
not gate_3207(n3283,n3282);
and gate_3208(n3284,pi38,n3283);
not gate_3209(n3285,n3284);
and gate_3210(n3286,n3268,n3285);
not gate_3211(n3287,n3286);
and gate_3212(n3288,n104,n3287);
and gate_3213(n3289,n81,n3288);
not gate_3214(n3290,n3289);
and gate_3215(n3291,n112,n148);
not gate_3216(n3292,n3291);
and gate_3217(n3293,pi06,n1105);
not gate_3218(n3294,n3293);
and gate_3219(n3295,n3292,n3294);
not gate_3220(n3296,n3295);
and gate_3221(n3297,pi38,n3296);
and gate_3222(n3298,pi34,n3297);
not gate_3223(n3299,n3298);
and gate_3224(n3300,n3290,n3299);
and gate_3225(n3301,n3254,n3300);
not gate_3226(n3302,n3301);
and gate_3227(n3303,n108,n3302);
not gate_3228(n3304,n3303);
and gate_3229(n3305,n129,n1722);
not gate_3230(n3306,n3305);
and gate_3231(n3307,n340,n3306);
not gate_3232(n3308,n3307);
and gate_3233(n3309,n129,n188);
not gate_3234(n3310,n3309);
and gate_3235(n3311,pi21,n3310);
not gate_3236(n3312,n3311);
and gate_3237(n3313,n1730,n3312);
and gate_3238(n3314,n3308,n3313);
not gate_3239(n3315,n3314);
and gate_3240(n3316,pi40,n3315);
not gate_3241(n3317,n3316);
and gate_3242(n3318,n1592,n3317);
not gate_3243(n3319,n3318);
and gate_3244(n3320,n692,n3319);
and gate_3245(n3321,pi15,n3320);
not gate_3246(n3322,n3321);
and gate_3247(n3323,n199,n625);
not gate_3248(n3324,n3323);
and gate_3249(n3325,n3322,n3324);
not gate_3250(n3326,n3325);
and gate_3251(n3327,n81,n3326);
not gate_3252(n3328,n3327);
and gate_3253(n3329,n110,n1905);
not gate_3254(n3330,n3329);
and gate_3255(n3331,n3328,n3330);
not gate_3256(n3332,n3331);
and gate_3257(n3333,n379,n3332);
not gate_3258(n3334,n3333);
and gate_3259(n3335,n3304,n3334);
not gate_3260(n3336,n3335);
and gate_3261(n3337,n109,n3336);
not gate_3262(n3338,n3337);
and gate_3263(n3339,n77,n535);
not gate_3264(n3340,n3339);
and gate_3265(n3341,pi01,n329);
not gate_3266(n3342,n3341);
and gate_3267(n3343,n3340,n3342);
not gate_3268(n3344,n3343);
and gate_3269(n3345,n2818,n3344);
and gate_3270(n3346,pi00,n3345);
not gate_3271(n3347,n3346);
and gate_3272(n3348,pi06,n1579);
not gate_3273(n3349,n3348);
and gate_3274(n3350,n615,n3349);
not gate_3275(n3351,n3350);
and gate_3276(n3352,pi40,n3351);
not gate_3277(n3353,n3352);
and gate_3278(n3354,n1598,n3353);
and gate_3279(n3355,n3347,n3354);
not gate_3280(n3356,n3355);
and gate_3281(n3357,pi35,n3356);
not gate_3282(n3358,n3357);
and gate_3283(n3359,n185,n1493);
not gate_3284(n3360,n3359);
and gate_3285(n3361,n184,n3360);
not gate_3286(n3362,n3361);
and gate_3287(n3363,n113,n3362);
not gate_3288(n3364,n3363);
and gate_3289(n3365,n720,n3122);
not gate_3290(n3366,n3365);
and gate_3291(n3367,n108,n3366);
not gate_3292(n3368,n3367);
and gate_3293(n3369,n220,n3368);
not gate_3294(n3370,n3369);
and gate_3295(n3371,n110,n3370);
not gate_3296(n3372,n3371);
and gate_3297(n3373,n3364,n3372);
and gate_3298(n3374,n3358,n3373);
not gate_3299(n3375,n3374);
and gate_3300(n3376,pi36,n3375);
not gate_3301(n3377,n3376);
and gate_3302(n3378,pi09,n104);
and gate_3303(n3379,n108,n181);
and gate_3304(n3380,n3378,n3379);
not gate_3305(n3381,n3380);
and gate_3306(n3382,n86,n87);
and gate_3307(n3383,n733,n3382);
not gate_3308(n3384,n3383);
and gate_3309(n3385,n3381,n3384);
not gate_3310(n3386,n3385);
and gate_3311(n3387,n85,n3386);
not gate_3312(n3388,n3387);
and gate_3313(n3389,n246,n3380);
not gate_3314(n3390,n3389);
and gate_3315(n3391,n87,n89);
not gate_3316(n3392,n3391);
and gate_3317(n3393,n2170,n3392);
not gate_3318(n3394,n3393);
and gate_3319(n3395,n733,n3394);
not gate_3320(n3396,n3395);
and gate_3321(n3397,n3390,n3396);
and gate_3322(n3398,n3388,n3397);
not gate_3323(n3399,n3398);
and gate_3324(n3400,n779,n3399);
and gate_3325(n3401,n81,n3400);
not gate_3326(n3402,n3401);
and gate_3327(n3403,n3377,n3402);
not gate_3328(n3404,n3403);
and gate_3329(n3405,n107,n3404);
not gate_3330(n3406,n3405);
and gate_3331(n3407,n3338,n3406);
not gate_3332(n3408,n3407);
and gate_3333(n3409,n105,n3408);
not gate_3334(n3410,n3409);
and gate_3335(n3411,n83,n3410);
not gate_3336(n3412,n3411);
and gate_3337(n3413,pi33,n3412);
not gate_3338(n3414,n3413);
and gate_3339(n3415,pi32,n106);
not gate_3340(n3416,n3415);
and gate_3341(n3417,n3414,n3416);
not gate_3342(po33,n3417);
and gate_3343(n3419,pi04,pi35);
not gate_3344(n3420,n3419);
and gate_3345(n3421,n108,n1423);
not gate_3346(n3422,n3421);
and gate_3347(n3423,n3420,n3422);
not gate_3348(n3424,n3423);
and gate_3349(n3425,n586,n3424);
and gate_3350(n3426,pi00,n3425);
not gate_3351(n3427,n3426);
and gate_3352(n3428,n1885,n2364);
not gate_3353(n3429,n3428);
and gate_3354(n3430,n3427,n3429);
not gate_3355(n3431,n3430);
and gate_3356(n3432,pi38,n3431);
not gate_3357(n3433,n3432);
and gate_3358(n3434,pi35,n1955);
not gate_3359(n3435,n3434);
and gate_3360(n3436,n113,n3435);
not gate_3361(n3437,n3436);
and gate_3362(n3438,pi06,n1461);
not gate_3363(n3439,n3438);
and gate_3364(n3440,n3437,n3439);
not gate_3365(n3441,n3440);
and gate_3366(n3442,n185,n3441);
not gate_3367(n3443,n3442);
and gate_3368(n3444,n3433,n3443);
not gate_3369(n3445,n3444);
and gate_3370(n3446,pi36,n3445);
not gate_3371(n3447,n3446);
and gate_3372(n3448,n197,n3236);
not gate_3373(n3449,n3448);
and gate_3374(n3450,n185,n3449);
and gate_3375(n3451,n170,n3450);
and gate_3376(n3452,n104,n3451);
not gate_3377(n3453,n3452);
and gate_3378(n3454,n3447,n3453);
not gate_3379(n3455,n3454);
and gate_3380(n3456,pi37,n3455);
not gate_3381(n3457,n3456);
and gate_3382(n3458,n109,n113);
not gate_3383(n3459,n3458);
and gate_3384(n3460,n1622,n3459);
not gate_3385(n3461,n3460);
and gate_3386(n3462,n76,n3461);
not gate_3387(n3463,n3462);
and gate_3388(n3464,n1892,n3463);
not gate_3389(n3465,n3464);
and gate_3390(n3466,pi05,n3465);
not gate_3391(n3467,n3466);
and gate_3392(n3468,n124,n2344);
not gate_3393(n3469,n3468);
and gate_3394(n3470,pi40,n3469);
not gate_3395(n3471,n3470);
and gate_3396(n3472,pi36,n3471);
not gate_3397(n3473,n3472);
and gate_3398(n3474,n113,n2222);
and gate_3399(n3475,n104,n3474);
not gate_3400(n3476,n3475);
and gate_3401(n3477,n510,n2221);
not gate_3402(n3478,n3477);
and gate_3403(n3479,pi31,n3478);
not gate_3404(n3480,n3479);
and gate_3405(n3481,pi40,n3480);
and gate_3406(n3482,n109,n3481);
and gate_3407(n3483,n263,n3482);
not gate_3408(n3484,n3483);
and gate_3409(n3485,n3476,n3484);
not gate_3410(n3486,n3485);
and gate_3411(n3487,pi09,n3486);
not gate_3412(n3488,n3487);
and gate_3413(n3489,n277,n3482);
not gate_3414(n3490,n3489);
and gate_3415(n3491,n3488,n3490);
and gate_3416(n3492,n3473,n3491);
not gate_3417(n3493,n3492);
and gate_3418(n3494,n108,n3493);
not gate_3419(n3495,n3494);
and gate_3420(n3496,pi36,n3438);
not gate_3421(n3497,n3496);
and gate_3422(n3498,n3495,n3497);
not gate_3423(n3499,n3498);
and gate_3424(n3500,n110,n3499);
not gate_3425(n3501,n3500);
and gate_3426(n3502,n3467,n3501);
not gate_3427(n3503,n3502);
and gate_3428(n3504,pi38,n3503);
not gate_3429(n3505,n3504);
and gate_3430(n3506,n198,n411);
not gate_3431(n3507,n3506);
and gate_3432(n3508,pi09,n89);
not gate_3433(n3509,n3508);
and gate_3434(n3510,n3507,n3509);
not gate_3435(n3511,n3510);
and gate_3436(n3512,n110,n3511);
and gate_3437(n3513,n104,n3512);
not gate_3438(n3514,n3513);
and gate_3439(n3515,n81,n3514);
not gate_3440(n3516,n3515);
and gate_3441(n3517,n109,n3516);
not gate_3442(n3518,n3517);
and gate_3443(n3519,n1443,n1645);
not gate_3444(n3520,n3519);
and gate_3445(n3521,n3518,n3520);
not gate_3446(n3522,n3521);
and gate_3447(n3523,n108,n3522);
not gate_3448(n3524,n3523);
and gate_3449(n3525,n109,n1173);
and gate_3450(n3526,n547,n3525);
not gate_3451(n3527,n3526);
and gate_3452(n3528,n3524,n3527);
and gate_3453(n3529,n3505,n3528);
not gate_3454(n3530,n3529);
and gate_3455(n3531,pi39,n3530);
not gate_3456(n3532,n3531);
and gate_3457(n3533,n496,n2555);
and gate_3458(n3534,n432,n3533);
not gate_3459(n3535,n3534);
and gate_3460(n3536,n108,n3535);
not gate_3461(n3537,n3536);
and gate_3462(n3538,pi37,n1462);
not gate_3463(n3539,n3538);
and gate_3464(n3540,n185,n3539);
not gate_3465(n3541,n3540);
and gate_3466(n3542,n3537,n3541);
not gate_3467(n3543,n3542);
and gate_3468(n3544,pi05,n3543);
not gate_3469(n3545,n3544);
and gate_3470(n3546,n108,n1173);
not gate_3471(n3547,n3546);
and gate_3472(n3548,n573,n3547);
not gate_3473(n3549,n3548);
and gate_3474(n3550,n198,n3549);
and gate_3475(n3551,n104,n3550);
not gate_3476(n3552,n3551);
and gate_3477(n3553,n526,n547);
not gate_3478(n3554,n3553);
and gate_3479(n3555,n3552,n3554);
and gate_3480(n3556,n3545,n3555);
not gate_3481(n3557,n3556);
and gate_3482(n3558,n109,n3557);
not gate_3483(n3559,n3558);
and gate_3484(n3560,n3532,n3559);
and gate_3485(n3561,n3457,n3560);
not gate_3486(n3562,n3561);
and gate_3487(n3563,n107,n3562);
not gate_3488(n3564,n3563);
and gate_3489(n3565,pi05,pi37);
and gate_3490(n3566,n400,n3565);
not gate_3491(n3567,n3566);
and gate_3492(n3568,pi34,n2344);
and gate_3493(n3569,n143,n3568);
not gate_3494(n3570,n3569);
and gate_3495(n3571,n1886,n3570);
not gate_3496(n3572,n3571);
and gate_3497(n3573,n2303,n3572);
not gate_3498(n3574,n3573);
and gate_3499(n3575,n3567,n3574);
not gate_3500(n3576,n3575);
and gate_3501(n3577,n111,n3576);
not gate_3502(n3578,n3577);
and gate_3503(n3579,n328,n2341);
not gate_3504(n3580,n3579);
and gate_3505(n3581,n535,n3580);
and gate_3506(n3582,pi34,n3581);
not gate_3507(n3583,n3582);
and gate_3508(n3584,n3578,n3583);
not gate_3509(n3585,n3584);
and gate_3510(n3586,n170,n3585);
not gate_3511(n3587,n3586);
and gate_3512(n3588,n3564,n3587);
not gate_3513(n3589,n3588);
and gate_3514(n3590,n105,n3589);
not gate_3515(n3591,n3590);
and gate_3516(n3592,n83,n3591);
not gate_3517(n3593,n3592);
and gate_3518(po34,pi33,n3593);
endmodule
