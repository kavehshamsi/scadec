
module c432_xrnd_32 ( G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, 
        G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, 
        G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, 
        G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, 
        G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, 
        G431gat, G432gat, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31 );
  input G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat,
         G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat,
         G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat,
         G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat,
         G108gat, G112gat, G115gat, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31;
  output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
  wire   n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327;

  NAND2_X1 U164 ( .A1(n163), .A2(n164), .ZN(G432gat) );
  NAND2_X1 U165 ( .A1(n165), .A2(n166), .ZN(n164) );
  MUX2_X1 U166 ( .A(n167), .B(n168), .S(keyinput18), .Z(n165) );
  NAND3_X1 U167 ( .A1(n169), .A2(n168), .A3(n170), .ZN(n167) );
  OR2_X1 U168 ( .A1(n171), .A2(n172), .ZN(n170) );
  NAND2_X1 U169 ( .A1(n173), .A2(n174), .ZN(n169) );
  XNOR2_X1 U170 ( .A(keyinput8), .B(n175), .ZN(n173) );
  NAND3_X1 U171 ( .A1(n163), .A2(n166), .A3(n176), .ZN(G431gat) );
  NAND3_X1 U172 ( .A1(n177), .A2(n168), .A3(n178), .ZN(n176) );
  NAND4_X1 U173 ( .A1(n179), .A2(n177), .A3(n163), .A4(n166), .ZN(G430gat) );
  XNOR2_X1 U174 ( .A(n180), .B(keyinput18), .ZN(n179) );
  NOR2_X1 U175 ( .A1(n181), .A2(n182), .ZN(G421gat) );
  NOR4_X1 U176 ( .A1(n183), .A2(n184), .A3(n185), .A4(n186), .ZN(n182) );
  NOR2_X1 U177 ( .A1(n187), .A2(n188), .ZN(n185) );
  AND2_X1 U178 ( .A1(G223gat), .A2(G1gat), .ZN(n184) );
  NOR2_X1 U179 ( .A1(n189), .A2(n190), .ZN(n183) );
  INV_X1 U180 ( .A(G370gat), .ZN(n189) );
  NOR4_X1 U181 ( .A1(n191), .A2(n178), .A3(n180), .A4(n172), .ZN(n181) );
  INV_X1 U182 ( .A(n177), .ZN(n172) );
  NAND4_X1 U183 ( .A1(G56gat), .A2(n192), .A3(n193), .A4(n194), .ZN(n177) );
  NAND2_X1 U184 ( .A1(n195), .A2(G329gat), .ZN(n194) );
  NAND2_X1 U185 ( .A1(G50gat), .A2(G223gat), .ZN(n193) );
  NAND2_X1 U186 ( .A1(G66gat), .A2(G370gat), .ZN(n192) );
  INV_X1 U187 ( .A(n168), .ZN(n180) );
  NAND4_X1 U188 ( .A1(G43gat), .A2(n196), .A3(n197), .A4(n198), .ZN(n168) );
  NAND2_X1 U189 ( .A1(G37gat), .A2(G223gat), .ZN(n198) );
  NAND2_X1 U190 ( .A1(G47gat), .A2(G329gat), .ZN(n197) );
  NAND2_X1 U191 ( .A1(G53gat), .A2(G370gat), .ZN(n196) );
  NAND2_X1 U192 ( .A1(n174), .A2(n171), .ZN(n178) );
  NAND4_X1 U193 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(n171) );
  XOR2_X1 U194 ( .A(n203), .B(keyinput24), .Z(n200) );
  NAND2_X1 U195 ( .A1(G73gat), .A2(G329gat), .ZN(n203) );
  XOR2_X1 U196 ( .A(n204), .B(keyinput1), .Z(n199) );
  NAND2_X1 U197 ( .A1(n205), .A2(G370gat), .ZN(n204) );
  NAND3_X1 U198 ( .A1(n206), .A2(n207), .A3(n208), .ZN(n174) );
  INV_X1 U199 ( .A(n209), .ZN(n208) );
  NAND2_X1 U200 ( .A1(n210), .A2(G370gat), .ZN(n207) );
  NAND2_X1 U201 ( .A1(G86gat), .A2(G329gat), .ZN(n206) );
  NAND4_X1 U202 ( .A1(n163), .A2(n166), .A3(n211), .A4(n175), .ZN(n191) );
  NAND4_X1 U203 ( .A1(n212), .A2(n213), .A3(n214), .A4(n215), .ZN(n175) );
  NAND2_X1 U204 ( .A1(n216), .A2(G370gat), .ZN(n214) );
  XOR2_X1 U205 ( .A(n217), .B(keyinput23), .Z(n212) );
  NAND2_X1 U206 ( .A1(G99gat), .A2(G329gat), .ZN(n217) );
  NAND4_X1 U207 ( .A1(G108gat), .A2(n218), .A3(n219), .A4(n220), .ZN(n211) );
  OR2_X1 U208 ( .A1(n221), .A2(n187), .ZN(n220) );
  NAND2_X1 U209 ( .A1(G115gat), .A2(G370gat), .ZN(n219) );
  NAND4_X1 U210 ( .A1(n222), .A2(n223), .A3(G30gat), .A4(n224), .ZN(n166) );
  NAND2_X1 U211 ( .A1(n225), .A2(G370gat), .ZN(n224) );
  XOR2_X1 U212 ( .A(n226), .B(keyinput29), .Z(n223) );
  NAND2_X1 U213 ( .A1(G34gat), .A2(G329gat), .ZN(n226) );
  XOR2_X1 U214 ( .A(n227), .B(n228), .Z(n222) );
  XOR2_X1 U215 ( .A(keyinput4), .B(keyinput28), .Z(n228) );
  NAND4_X1 U216 ( .A1(G17gat), .A2(n229), .A3(n230), .A4(n231), .ZN(n163) );
  NAND2_X1 U217 ( .A1(G21gat), .A2(G329gat), .ZN(n230) );
  NAND2_X1 U218 ( .A1(G27gat), .A2(G370gat), .ZN(n229) );
  NAND4_X1 U219 ( .A1(n232), .A2(n233), .A3(n234), .A4(n235), .ZN(G370gat) );
  NAND4_X1 U220 ( .A1(n236), .A2(n237), .A3(n238), .A4(n239), .ZN(n235) );
  INV_X1 U221 ( .A(G53gat), .ZN(n239) );
  XNOR2_X1 U222 ( .A(n240), .B(n241), .ZN(n236) );
  XNOR2_X1 U223 ( .A(n242), .B(keyinput22), .ZN(n241) );
  NOR2_X1 U224 ( .A1(n243), .A2(n244), .ZN(n234) );
  NOR4_X1 U225 ( .A1(n245), .A2(n246), .A3(n247), .A4(n205), .ZN(n244) );
  XOR2_X1 U226 ( .A(keyinput25), .B(G79gat), .Z(n205) );
  XNOR2_X1 U227 ( .A(n240), .B(n248), .ZN(n247) );
  NOR3_X1 U228 ( .A1(n210), .A2(n249), .A3(n209), .ZN(n243) );
  XNOR2_X1 U229 ( .A(n240), .B(n250), .ZN(n249) );
  XOR2_X1 U230 ( .A(keyinput12), .B(G92gat), .Z(n210) );
  XOR2_X1 U231 ( .A(n251), .B(keyinput0), .Z(n233) );
  NAND3_X1 U232 ( .A1(n252), .A2(n231), .A3(n253), .ZN(n251) );
  XOR2_X1 U233 ( .A(keyinput20), .B(n254), .Z(n253) );
  NOR2_X1 U234 ( .A1(G27gat), .A2(n255), .ZN(n254) );
  XNOR2_X1 U235 ( .A(n256), .B(n257), .ZN(n252) );
  MUX2_X1 U236 ( .A(n258), .B(n259), .S(n257), .Z(n232) );
  INV_X1 U237 ( .A(n240), .ZN(n257) );
  XOR2_X1 U238 ( .A(n187), .B(keyinput14), .Z(n240) );
  NOR4_X1 U239 ( .A1(n260), .A2(n261), .A3(n262), .A4(n263), .ZN(n259) );
  NOR2_X1 U240 ( .A1(n264), .A2(n265), .ZN(n263) );
  INV_X1 U241 ( .A(n266), .ZN(n265) );
  NOR2_X1 U242 ( .A1(n267), .A2(n268), .ZN(n262) );
  NAND2_X1 U243 ( .A1(n269), .A2(n270), .ZN(n261) );
  NAND2_X1 U244 ( .A1(n271), .A2(n190), .ZN(n270) );
  NAND2_X1 U245 ( .A1(n272), .A2(n273), .ZN(n269) );
  INV_X1 U246 ( .A(n216), .ZN(n273) );
  NOR2_X1 U247 ( .A1(n274), .A2(n275), .ZN(n260) );
  INV_X1 U248 ( .A(n276), .ZN(n274) );
  NOR3_X1 U249 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n258) );
  NOR2_X1 U250 ( .A1(n266), .A2(n264), .ZN(n279) );
  XOR2_X1 U251 ( .A(n280), .B(keyinput3), .Z(n264) );
  NAND3_X1 U252 ( .A1(n281), .A2(n227), .A3(n282), .ZN(n280) );
  XOR2_X1 U253 ( .A(keyinput2), .B(n283), .Z(n282) );
  NOR2_X1 U254 ( .A1(n284), .A2(n225), .ZN(n283) );
  XOR2_X1 U255 ( .A(keyinput19), .B(G40gat), .Z(n225) );
  NAND2_X1 U256 ( .A1(G223gat), .A2(n284), .ZN(n281) );
  NOR2_X1 U257 ( .A1(n285), .A2(n267), .ZN(n278) );
  XOR2_X1 U258 ( .A(n286), .B(keyinput15), .Z(n267) );
  NAND3_X1 U259 ( .A1(n218), .A2(n287), .A3(G108gat), .ZN(n286) );
  INV_X1 U260 ( .A(G115gat), .ZN(n287) );
  NAND3_X1 U261 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n277) );
  NAND2_X1 U262 ( .A1(n275), .A2(n276), .ZN(n290) );
  XNOR2_X1 U263 ( .A(n291), .B(keyinput17), .ZN(n276) );
  NAND2_X1 U264 ( .A1(n292), .A2(n293), .ZN(n291) );
  XOR2_X1 U265 ( .A(keyinput11), .B(n294), .Z(n292) );
  NOR2_X1 U266 ( .A1(G66gat), .A2(n295), .ZN(n294) );
  XNOR2_X1 U267 ( .A(n296), .B(keyinput10), .ZN(n275) );
  NAND3_X1 U268 ( .A1(n297), .A2(n298), .A3(n190), .ZN(n289) );
  XNOR2_X1 U269 ( .A(keyinput7), .B(G14gat), .ZN(n190) );
  OR3_X1 U270 ( .A1(n299), .A2(n272), .A3(n216), .ZN(n288) );
  XOR2_X1 U271 ( .A(keyinput16), .B(G105gat), .Z(n216) );
  INV_X1 U272 ( .A(n187), .ZN(G329gat) );
  NOR4_X1 U273 ( .A1(n250), .A2(n248), .A3(n300), .A4(n301), .ZN(n187) );
  OR4_X1 U274 ( .A1(n272), .A2(n285), .A3(n296), .A4(n242), .ZN(n301) );
  AND3_X1 U275 ( .A1(n238), .A2(n302), .A3(n237), .ZN(n242) );
  XNOR2_X1 U276 ( .A(n303), .B(G43gat), .ZN(n237) );
  XNOR2_X1 U277 ( .A(keyinput9), .B(keyinput30), .ZN(n303) );
  INV_X1 U278 ( .A(G47gat), .ZN(n302) );
  NAND2_X1 U279 ( .A1(G223gat), .A2(n304), .ZN(n238) );
  NAND2_X1 U280 ( .A1(G43gat), .A2(n305), .ZN(n304) );
  NOR3_X1 U281 ( .A1(n295), .A2(n306), .A3(n195), .ZN(n296) );
  XOR2_X1 U282 ( .A(keyinput27), .B(G60gat), .Z(n195) );
  INV_X1 U283 ( .A(n293), .ZN(n306) );
  XNOR2_X1 U284 ( .A(n307), .B(n308), .ZN(n293) );
  XOR2_X1 U285 ( .A(G223gat), .B(keyinput6), .Z(n307) );
  INV_X1 U286 ( .A(n268), .ZN(n285) );
  NAND3_X1 U287 ( .A1(G108gat), .A2(n218), .A3(n221), .ZN(n268) );
  XNOR2_X1 U288 ( .A(keyinput21), .B(G112gat), .ZN(n221) );
  NAND2_X1 U289 ( .A1(G102gat), .A2(G223gat), .ZN(n218) );
  NOR2_X1 U290 ( .A1(n299), .A2(G99gat), .ZN(n272) );
  NAND2_X1 U291 ( .A1(n213), .A2(n215), .ZN(n299) );
  NAND2_X1 U292 ( .A1(G89gat), .A2(G223gat), .ZN(n215) );
  OR3_X1 U293 ( .A1(n256), .A2(n266), .A3(n271), .ZN(n300) );
  INV_X1 U294 ( .A(n298), .ZN(n271) );
  NAND2_X1 U295 ( .A1(n297), .A2(n188), .ZN(n298) );
  INV_X1 U296 ( .A(G8gat), .ZN(n188) );
  AND2_X1 U297 ( .A1(G4gat), .A2(n309), .ZN(n297) );
  NAND2_X1 U298 ( .A1(G1gat), .A2(G223gat), .ZN(n309) );
  NOR3_X1 U299 ( .A1(n310), .A2(G34gat), .A3(n284), .ZN(n266) );
  INV_X1 U300 ( .A(n227), .ZN(n310) );
  NAND2_X1 U301 ( .A1(G24gat), .A2(G223gat), .ZN(n227) );
  NOR3_X1 U302 ( .A1(n311), .A2(G21gat), .A3(n255), .ZN(n256) );
  INV_X1 U303 ( .A(G17gat), .ZN(n255) );
  INV_X1 U304 ( .A(n231), .ZN(n311) );
  NAND2_X1 U305 ( .A1(G223gat), .A2(n312), .ZN(n231) );
  NOR3_X1 U306 ( .A1(n245), .A2(G73gat), .A3(n246), .ZN(n248) );
  INV_X1 U307 ( .A(n201), .ZN(n246) );
  INV_X1 U308 ( .A(n202), .ZN(n245) );
  NAND2_X1 U309 ( .A1(G223gat), .A2(n313), .ZN(n202) );
  NOR2_X1 U310 ( .A1(n209), .A2(G86gat), .ZN(n250) );
  NAND2_X1 U311 ( .A1(G82gat), .A2(n314), .ZN(n209) );
  NAND2_X1 U312 ( .A1(G76gat), .A2(G223gat), .ZN(n314) );
  NAND4_X1 U313 ( .A1(n315), .A2(n316), .A3(n317), .A4(n318), .ZN(G223gat) );
  NOR4_X1 U314 ( .A1(n319), .A2(n320), .A3(n308), .A4(n321), .ZN(n318) );
  NOR2_X1 U315 ( .A1(G76gat), .A2(n322), .ZN(n321) );
  INV_X1 U316 ( .A(G82gat), .ZN(n322) );
  NOR2_X1 U317 ( .A1(G50gat), .A2(n295), .ZN(n308) );
  INV_X1 U318 ( .A(G56gat), .ZN(n295) );
  AND2_X1 U319 ( .A1(n305), .A2(G43gat), .ZN(n320) );
  INV_X1 U320 ( .A(G37gat), .ZN(n305) );
  NOR2_X1 U321 ( .A1(G24gat), .A2(n284), .ZN(n319) );
  INV_X1 U322 ( .A(G30gat), .ZN(n284) );
  AND3_X1 U323 ( .A1(n323), .A2(n313), .A3(n312), .ZN(n317) );
  NAND2_X1 U324 ( .A1(n324), .A2(G17gat), .ZN(n312) );
  XNOR2_X1 U325 ( .A(keyinput13), .B(G11gat), .ZN(n324) );
  NAND2_X1 U326 ( .A1(n325), .A2(n201), .ZN(n313) );
  XOR2_X1 U327 ( .A(keyinput26), .B(G69gat), .Z(n201) );
  XNOR2_X1 U328 ( .A(keyinput31), .B(G63gat), .ZN(n325) );
  NAND2_X1 U329 ( .A1(n326), .A2(n213), .ZN(n323) );
  XOR2_X1 U330 ( .A(keyinput5), .B(G95gat), .Z(n213) );
  INV_X1 U331 ( .A(G89gat), .ZN(n326) );
  NAND2_X1 U332 ( .A1(G108gat), .A2(n327), .ZN(n316) );
  INV_X1 U333 ( .A(G102gat), .ZN(n327) );
  OR2_X1 U334 ( .A1(n186), .A2(G1gat), .ZN(n315) );
  INV_X1 U335 ( .A(G4gat), .ZN(n186) );
endmodule

