module c432 ( G432gat, G431gat, G430gat, G421gat, G370gat, G329gat, G223gat, 
        G115gat, G112gat, G108gat, G105gat, G102gat, G99gat, G95gat, G92gat, 
        G89gat, G86gat, G82gat, G79gat, G76gat, G73gat, G30gat, G27gat, G24gat, 
        G21gat, G17gat, G14gat, G11gat, G8gat, G4gat, G1gat, G34gat, G37gat, 
        G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, 
        G69gat );
  input G115gat, G112gat, G108gat, G105gat, G102gat, G99gat, G95gat, G92gat,
         G89gat, G86gat, G82gat, G79gat, G76gat, G73gat, G30gat, G27gat,
         G24gat, G21gat, G17gat, G14gat, G11gat, G8gat, G4gat, G1gat, G34gat,
         G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat,
         G63gat, G66gat, G69gat;
  output G432gat, G431gat, G430gat, G421gat, G370gat, G329gat, G223gat;
  wire   n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179;

  INV_X1 U94 ( .A(G1gat), .ZN(n97) );
  INV_X1 U95 ( .A(G43gat), .ZN(n114) );
  NOR2_X1 U96 ( .A1(G37gat), .A2(n114), .ZN(n151) );
  AOI21_X1 U97 ( .B1(G4gat), .B2(n97), .A(n151), .ZN(n95) );
  INV_X1 U98 ( .A(G102gat), .ZN(n101) );
  INV_X1 U99 ( .A(G30gat), .ZN(n146) );
  NOR2_X1 U100 ( .A1(G24gat), .A2(n146), .ZN(n124) );
  INV_X1 U101 ( .A(G56gat), .ZN(n111) );
  NOR2_X1 U102 ( .A1(G50gat), .A2(n111), .ZN(n153) );
  AOI211_X1 U103 ( .C1(G108gat), .C2(n101), .A(n124), .B(n153), .ZN(n94) );
  INV_X1 U104 ( .A(G95gat), .ZN(n118) );
  NOR2_X1 U105 ( .A1(G89gat), .A2(n118), .ZN(n96) );
  INV_X1 U106 ( .A(G17gat), .ZN(n98) );
  NOR2_X1 U107 ( .A1(G11gat), .A2(n98), .ZN(n148) );
  INV_X1 U108 ( .A(G82gat), .ZN(n110) );
  NOR2_X1 U109 ( .A1(G76gat), .A2(n110), .ZN(n162) );
  INV_X1 U110 ( .A(G69gat), .ZN(n115) );
  NOR2_X1 U111 ( .A1(G63gat), .A2(n115), .ZN(n102) );
  NOR4_X1 U112 ( .A1(n96), .A2(n148), .A3(n162), .A4(n102), .ZN(n93) );
  NAND3_X1 U113 ( .A1(n95), .A2(n94), .A3(n93), .ZN(G223gat) );
  INV_X1 U114 ( .A(G223gat), .ZN(n161) );
  AOI21_X1 U115 ( .B1(G95gat), .B2(n161), .A(n96), .ZN(n157) );
  OAI21_X1 U116 ( .B1(n161), .B2(n97), .A(G4gat), .ZN(n154) );
  NOR2_X1 U117 ( .A1(G8gat), .A2(n154), .ZN(n120) );
  AOI211_X1 U118 ( .C1(G11gat), .C2(G223gat), .A(G21gat), .B(n98), .ZN(n119)
         );
  INV_X1 U119 ( .A(G60gat), .ZN(n112) );
  OAI22_X1 U120 ( .A1(G73gat), .A2(n115), .B1(G47gat), .B2(n114), .ZN(n100) );
  OAI22_X1 U121 ( .A1(G86gat), .A2(n110), .B1(G34gat), .B2(n146), .ZN(n99) );
  AOI211_X1 U122 ( .C1(G56gat), .C2(n112), .A(n100), .B(n99), .ZN(n107) );
  INV_X1 U123 ( .A(G86gat), .ZN(n113) );
  AOI22_X1 U124 ( .A1(n162), .A2(n113), .B1(n153), .B2(n112), .ZN(n106) );
  INV_X1 U125 ( .A(G47gat), .ZN(n117) );
  OAI21_X1 U126 ( .B1(n161), .B2(n101), .A(G108gat), .ZN(n165) );
  NOR2_X1 U127 ( .A1(G112gat), .A2(n165), .ZN(n125) );
  INV_X1 U128 ( .A(n124), .ZN(n103) );
  INV_X1 U129 ( .A(n102), .ZN(n158) );
  OAI22_X1 U130 ( .A1(G34gat), .A2(n103), .B1(G73gat), .B2(n158), .ZN(n104) );
  AOI211_X1 U131 ( .C1(n151), .C2(n117), .A(n125), .B(n104), .ZN(n105) );
  OAI211_X1 U132 ( .C1(n107), .C2(G223gat), .A(n106), .B(n105), .ZN(n108) );
  NOR3_X1 U133 ( .A1(n120), .A2(n119), .A3(n108), .ZN(n109) );
  OAI21_X1 U134 ( .B1(G99gat), .B2(n157), .A(n109), .ZN(G329gat) );
  AOI211_X1 U135 ( .C1(G76gat), .C2(G223gat), .A(G92gat), .B(n110), .ZN(n131)
         );
  AOI211_X1 U136 ( .C1(G50gat), .C2(G223gat), .A(G66gat), .B(n111), .ZN(n130)
         );
  AOI22_X1 U137 ( .A1(n131), .A2(n113), .B1(n130), .B2(n112), .ZN(n143) );
  AOI211_X1 U138 ( .C1(G37gat), .C2(G223gat), .A(G53gat), .B(n114), .ZN(n132)
         );
  AOI211_X1 U139 ( .C1(G63gat), .C2(G223gat), .A(G79gat), .B(n115), .ZN(n133)
         );
  INV_X1 U140 ( .A(G73gat), .ZN(n116) );
  AOI22_X1 U141 ( .A1(n132), .A2(n117), .B1(n133), .B2(n116), .ZN(n142) );
  AOI211_X1 U142 ( .C1(G89gat), .C2(G223gat), .A(G105gat), .B(n118), .ZN(n129)
         );
  NAND2_X1 U143 ( .A1(G99gat), .A2(G329gat), .ZN(n155) );
  INV_X1 U144 ( .A(n119), .ZN(n122) );
  INV_X1 U145 ( .A(n120), .ZN(n121) );
  OAI22_X1 U146 ( .A1(G27gat), .A2(n122), .B1(G14gat), .B2(n121), .ZN(n128) );
  INV_X1 U147 ( .A(G40gat), .ZN(n123) );
  OAI211_X1 U148 ( .C1(n124), .C2(n161), .A(G30gat), .B(n123), .ZN(n134) );
  INV_X1 U149 ( .A(n125), .ZN(n126) );
  OAI22_X1 U150 ( .A1(G34gat), .A2(n134), .B1(G115gat), .B2(n126), .ZN(n127)
         );
  AOI211_X1 U151 ( .C1(n129), .C2(n155), .A(n128), .B(n127), .ZN(n141) );
  OAI22_X1 U152 ( .A1(G14gat), .A2(n154), .B1(G115gat), .B2(n165), .ZN(n139)
         );
  OAI21_X1 U153 ( .B1(n148), .B2(n161), .A(G17gat), .ZN(n136) );
  NOR4_X1 U154 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(n135) );
  OAI211_X1 U155 ( .C1(G27gat), .C2(n136), .A(n135), .B(n134), .ZN(n138) );
  INV_X1 U156 ( .A(G329gat), .ZN(n137) );
  OAI21_X1 U157 ( .B1(n139), .B2(n138), .A(n137), .ZN(n140) );
  NAND4_X1 U158 ( .A1(n143), .A2(n142), .A3(n141), .A4(n140), .ZN(G370gat) );
  AOI22_X1 U159 ( .A1(G329gat), .A2(G34gat), .B1(G370gat), .B2(G40gat), .ZN(
        n144) );
  INV_X1 U160 ( .A(n144), .ZN(n145) );
  AOI211_X1 U161 ( .C1(G24gat), .C2(G223gat), .A(n146), .B(n145), .ZN(n179) );
  AOI22_X1 U162 ( .A1(G21gat), .A2(G329gat), .B1(G27gat), .B2(G370gat), .ZN(
        n147) );
  OAI211_X1 U163 ( .C1(n148), .C2(n161), .A(G17gat), .B(n147), .ZN(n176) );
  INV_X1 U164 ( .A(n176), .ZN(n149) );
  NOR2_X1 U165 ( .A1(n179), .A2(n149), .ZN(n169) );
  AOI22_X1 U166 ( .A1(G47gat), .A2(G329gat), .B1(G53gat), .B2(G370gat), .ZN(
        n150) );
  OAI211_X1 U167 ( .C1(n151), .C2(n161), .A(G43gat), .B(n150), .ZN(n177) );
  AOI22_X1 U168 ( .A1(G60gat), .A2(G329gat), .B1(G66gat), .B2(G370gat), .ZN(
        n152) );
  OAI211_X1 U169 ( .C1(n153), .C2(n161), .A(G56gat), .B(n152), .ZN(n172) );
  NAND3_X1 U170 ( .A1(n169), .A2(n177), .A3(n172), .ZN(G430gat) );
  INV_X1 U171 ( .A(n154), .ZN(n168) );
  AOI22_X1 U172 ( .A1(G8gat), .A2(G329gat), .B1(G14gat), .B2(G370gat), .ZN(
        n167) );
  INV_X1 U173 ( .A(n155), .ZN(n156) );
  AOI211_X1 U174 ( .C1(G105gat), .C2(G370gat), .A(n157), .B(n156), .ZN(n175)
         );
  NAND2_X1 U175 ( .A1(G69gat), .A2(n161), .ZN(n159) );
  AOI222_X1 U176 ( .A1(n159), .A2(n158), .B1(G329gat), .B2(G73gat), .C1(
        G370gat), .C2(G79gat), .ZN(n173) );
  AOI22_X1 U177 ( .A1(G86gat), .A2(G329gat), .B1(G92gat), .B2(G370gat), .ZN(
        n160) );
  OAI211_X1 U178 ( .C1(n162), .C2(n161), .A(G82gat), .B(n160), .ZN(n174) );
  INV_X1 U179 ( .A(n174), .ZN(n163) );
  NOR2_X1 U180 ( .A1(n173), .A2(n163), .ZN(n171) );
  INV_X1 U181 ( .A(n171), .ZN(n164) );
  NOR3_X1 U182 ( .A1(n175), .A2(n164), .A3(G430gat), .ZN(n166) );
  AOI22_X1 U183 ( .A1(n168), .A2(n167), .B1(n166), .B2(n165), .ZN(G421gat) );
  NAND2_X1 U184 ( .A1(n177), .A2(n172), .ZN(n170) );
  OAI21_X1 U185 ( .B1(n171), .B2(n170), .A(n169), .ZN(G431gat) );
  AOI22_X1 U186 ( .A1(n175), .A2(n174), .B1(n173), .B2(n172), .ZN(n178) );
  OAI221_X1 U187 ( .B1(n179), .B2(n178), .C1(n179), .C2(n177), .A(n176), .ZN(
        G432gat) );
endmodule

