// Verilog File 
module c3540 (G1,G13,G20,G33,G41,G45,G50,G58,G68,
G77,G87,G97,G107,G116,G124,G125,G128,G132,G137,
G143,G150,G159,G169,G179,G190,G200,G213,G222,G223,
G226,G232,G238,G244,G250,G257,G264,G270,G274,G283,
G294,G303,G311,G317,G322,G326,G329,G330,G343,G1698,
G2897,G353,G355,G361,G358,G351,G372,G369,G399,G364,
G396,G384,G367,G387,G393,G390,G378,G375,G381,G407,
G409,G405,G402);

input G1,G13,G20,G33,G41,G45,G50,G58,G68,
G77,G87,G97,G107,G116,G124,G125,G128,G132,G137,
G143,G150,G159,G169,G179,G190,G200,G213,G222,G223,
G226,G232,G238,G244,G250,G257,G264,G270,G274,G283,
G294,G303,G311,G317,G322,G326,G329,G330,G343,G1698,
G2897;

output G353,G355,G361,G358,G351,G372,G369,G399,G364,
G396,G384,G367,G387,G393,G390,G378,G375,G381,G407,
G409,G405,G402;

wire G432,G442,G447,G456,G460,G463,G467,G476,G479,
G483,G492,G501,G504,G513,G517,G526,G530,G540,G587,
G704,G707,G714,G717,G724,G731,G732,G736,G741,G758,
G776,G780,G788,G791,G798,G799,G802,G826,G828,G831,
G833,G836,G839,G842,G845,G848,G851,G890,G898,G907,
G1032,G1035,G1048,G1049,G1050,G1051,G1540,G1699,G1826,G1827,
G1828,G2051,G2478,G2865,G2868,G2931,G2934,G2939,G2942,G2947,
G2950,G2957,G2960,G3007,G3079,G3087,G3095,G3103,G3419,G588,
G759,G1541,G1772,G1829,G1834,G2052,G625,G545,G546,G547,
G548,G549,G550,G551,G552,G2937,G2938,G2945,G2946,G621,
G626,G635,G636,G3085,G3101,G657,G675,G721,G784,G794,
G807,G816,G823,G860,G861,G864,G893,G896,G897,G3093,
G905,G906,G3109,G973,G980,G987,G994,G1001,G1008,G1015,
G1022,G1038,G1043,G1054,G1057,G1512,G1681,G1717,G1724,G1731,
G1738,G1745,G1752,G1759,G1766,G1773,G1790,G1808,G2278,G2481,
G3425,G2871,G2874,G2953,G2954,G2963,G2964,G3010,G3013,G3017,
G3020,G3027,G3030,G3037,G3040,G3082,G3090,G3098,G3106,G352,
G553,G554,G555,G556,G560,G561,G650,G956,G974,G975,
G976,G981,G982,G988,G989,G990,G995,G996,G997,G1002,
G1003,G1004,G1009,G1010,G1016,G1017,G1018,G1023,G1024,G1025,
G1720,G1727,G1734,G1741,G1748,G1755,G1762,G1769,G1791,G1809,
G1851,G1901,G1952,G2002,G2057,G2109,G2162,G2214,G2955,G2956,
G2965,G2966,G354,G557,G562,G586,G630,G634,G639,G642,
G3086,G644,G646,G3102,G654,G660,G678,G804,G806,G855,
G867,G903,G3094,G912,G3110,G915,G927,G941,G977,G978,
G984,G985,G991,G992,G998,G999,G1005,G1006,G1012,G1013,
G1019,G1020,G1026,G1027,G1060,G1063,G1066,G1069,G1527,G1530,
G1542,G1563,G1572,G1581,G1585,G1589,G1593,G1597,G1601,G1605,
G1716,G1718,G1723,G1725,G1730,G1732,G1737,G1739,G1744,G1746,
G1751,G1753,G1758,G1760,G1765,G1767,G1852,G1856,G1870,G1902,
G1906,G1920,G1953,G1957,G1971,G2003,G2007,G2021,G2058,G2062,
G2076,G2110,G2114,G2128,G2163,G2167,G2181,G2215,G2219,G2233,
G2285,G2288,G2289,G2293,G2298,G2302,G2877,G2983,G2986,G3014,
G3015,G3023,G3024,G3033,G3034,G3043,G3044,G643,G647,G680,
G904,G913,G920,G979,G993,G1000,G1007,G1021,G1028,G1719,
G1721,G1726,G1728,G1733,G1735,G1740,G1742,G1747,G1749,G1754,
G1756,G1761,G1763,G1768,G1770,G1794,G1799,G1812,G1817,G1859,
G1909,G1960,G2010,G2065,G2117,G2170,G2222,G2678,G2697,G2716,
G2733,G2751,G2768,G2785,G2802,G3016,G3025,G3026,G3035,G3036,
G3045,G3046,G2989,G2990,G610,G613,G616,G640,G648,G655,
G665,G668,G671,G683,G685,G688,G694,G696,G699,G870,
G887,G901,G910,G914,G916,G942,G943,G1072,G1084,G1096,
G1108,G1120,G1132,G1144,G1156,G1533,G1534,G1535,G1545,G1554,
G1610,G1619,G1628,G1637,G1646,G1655,G1664,G1673,G1722,G1729,
G1736,G1743,G1750,G1757,G1764,G1771,G1853,G1954,G2004,G2059,
G2164,G2216,G2485,G2900,G2903,G2967,G2970,G2975,G2978,G3047,
G3050,G3055,G3058,G574,G575,G617,G641,G649,G662,G672,
G690,G691,G701,G702,G902,G911,G917,G923,G1538,G1871,
G1872,G1873,G1921,G1922,G1923,G1972,G1973,G1974,G2022,G2023,
G2024,G2077,G2078,G2079,G2129,G2130,G2131,G2182,G2183,G2184,
G2234,G2235,G2236,G2973,G2974,G2981,G2982,G576,G3053,G3054,
G3061,G3062,G645,G926,G928,G947,G983,G1011,G1075,G1087,
G1099,G1111,G1123,G1135,G1147,G1159,G1168,G1177,G1186,G1195,
G1204,G1213,G1222,G1231,G1609,G1611,G1618,G1620,G1627,G1629,
G1636,G1638,G1645,G1647,G1654,G1656,G1663,G1665,G1672,G1674,
G1862,G1866,G1874,G1924,G1963,G1967,G1975,G2013,G2017,G2025,
G2068,G2072,G2080,G2132,G2173,G2177,G2185,G2225,G2229,G2237,
G2488,G2679,G2680,G2698,G2699,G2717,G2718,G2734,G2735,G2752,
G2753,G2769,G2770,G2786,G2787,G2803,G2804,G359,G1029,G565,
G566,G569,G570,G589,G590,G595,G596,G929,G938,G944,
G986,G1014,G1616,G1625,G1634,G1643,G360,G567,G571,G579,
G591,G597,G614,G1240,G1241,G1242,G1243,G1244,G1245,G1246,
G1247,G1257,G1258,G1259,G1260,G1261,G1262,G1263,G1264,G1274,
G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1291,G1292,G1293,
G1294,G1295,G1296,G1297,G1298,G1308,G1309,G1310,G1311,G1312,
G1313,G1314,G1315,G1325,G1326,G1327,G1328,G1329,G1330,G1331,
G1332,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1359,
G1360,G1361,G1362,G1363,G1364,G1365,G1366,G1376,G1377,G1378,
G1379,G1380,G1381,G1382,G1383,G1393,G1394,G1395,G1396,G1397,
G1398,G1399,G1400,G1410,G1411,G1412,G1413,G1414,G1415,G1416,
G1417,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1444,
G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1461,G1462,G1463,
G1464,G1465,G1466,G1467,G1468,G1478,G1479,G1480,G1481,G1482,
G1483,G1484,G1485,G1495,G1496,G1497,G1498,G1499,G1500,G1501,
G1502,G1877,G1880,G1891,G1903,G1927,G1930,G1978,G1981,G1992,
G2028,G2031,G2042,G2085,G2088,G2099,G2111,G2137,G2140,G2190,
G2193,G2204,G2242,G2245,G2256,G2320,G2341,G2354,G2367,G2383,
G2391,G2474,G2475,G2476,G2477,G2482,G568,G618,G1248,G1249,
G1250,G1251,G1252,G1253,G1254,G1255,G1265,G1266,G1267,G1268,
G1269,G1270,G1271,G1272,G1282,G1283,G1284,G1285,G1286,G1287,
G1288,G1289,G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,
G1316,G1317,G1318,G1319,G1320,G1321,G1322,G1323,G1333,G1334,
G1335,G1336,G1337,G1338,G1339,G1340,G1350,G1351,G1352,G1353,
G1354,G1355,G1356,G1357,G1367,G1368,G1369,G1370,G1371,G1372,
G1373,G1374,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,
G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408,G1418,G1419,
G1420,G1421,G1422,G1423,G1424,G1425,G1435,G1436,G1437,G1438,
G1439,G1440,G1441,G1442,G1452,G1453,G1454,G1455,G1456,G1457,
G1458,G1459,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,
G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,G1503,G1504,
G1505,G1506,G1507,G1508,G1509,G1510,G2483,G600,G661,G669,
G679,G1256,G1273,G1290,G1307,G1324,G1341,G1358,G1375,G1392,
G1409,G1426,G1443,G1460,G1477,G1494,G1511,G1652,G1883,G1886,
G1889,G1890,G1912,G1916,G1984,G1987,G1990,G1991,G2034,G2037,
G2040,G2041,G2091,G2094,G2097,G2098,G2120,G2124,G2196,G2199,
G2202,G2203,G2248,G2251,G2254,G2255,G2484,G2991,G2994,G2999,
G3002,G3063,G3071,G3124,G3134,G3158,G3166,G3174,G3182,G3190,
G3200,G3224,G3232,G3240,G3248,G663,G673,G681,G1536,G1537,
G1582,G1583,G1586,G1587,G1590,G1591,G1594,G1595,G1598,G1599,
G1602,G1603,G1606,G1607,G1894,G1997,G2047,G2102,G2209,G2261,
G2489,G3005,G3006,G3077,G3069,G2997,G2998,G689,G700,G1539,
G1584,G1588,G1592,G1596,G1600,G1604,G1608,G1661,G1892,G1893,
G1933,G1936,G1939,G1940,G1941,G1993,G1996,G2043,G2046,G2100,
G2101,G2143,G2146,G2149,G2150,G2151,G2205,G2208,G2257,G2260,
G3138,G2328,G3162,G3170,G3178,G3186,G3204,G2375,G3236,G3244,
G3252,G3228,G3066,G3074,G3128,G3194,G619,G620,G582,G583,
G692,G703,G1612,G1621,G1630,G1639,G1648,G1657,G1666,G1675,
G1895,G1946,G1998,G2048,G2103,G2156,G2210,G2262,G2271,G2311,
G356,G357,G603,G3078,G606,G3070,G1670,G1679,G1942,G1945,
G2152,G2155,G2445,G2448,G2455,G2458,G3142,G3150,G3208,G3216,
G604,G607,G1947,G2157,G2317,G2338,G2351,G2364,G2380,G2388,
G605,G608,G2272,G2312,G3146,G3154,G3220,G3212,G2444,G2451,
G2454,G2461,G2530,G3323,G349,G350,G2265,G2273,G2274,G2309,
G2313,G2314,G2325,G2372,G2523,G2533,G3121,G3131,G3155,G3163,
G3171,G3179,G3187,G3197,G3221,G3229,G3237,G3245,G2275,G2315,
G3329,G2324,G2350,G2363,G2371,G2387,G2400,G2268,G3137,G3161,
G2345,G3169,G3177,G2358,G3185,G3203,G3235,G3243,G2395,G3251,
G3227,G2432,G2490,G3127,G3130,G3139,G3147,G3193,G3196,G3205,
G3213,G2307,G2308,G2323,G2349,G2362,G2370,G2386,G2399,G2344,
G2357,G2394,G2431,G2464,G2491,G3129,G3195,G368,G1615,G2337,
G1633,G1642,G1651,G2379,G1669,G1678,G3145,G2332,G3153,G2346,
G2359,G3219,G2396,G3211,G2425,G2433,G3272,G3308,G1613,G2336,
G1631,G1640,G1649,G2378,G1667,G1676,G2331,G2424,G2467,G2495,
G3295,G3374,G1614,G1624,G1632,G1641,G1650,G1660,G1668,G1677,
G2333,G2406,G2409,G2415,G2419,G2426,G2439,G2518,G3276,G3312,
G2612,G3326,G1617,G1622,G1635,G1644,G1653,G1658,G1671,G1680,
G2500,G2505,G2519,G3378,G2642,G2645,G3301,G1623,G1659,G2401,
G2501,G2511,G2512,G2513,G2514,G2517,G2531,G2532,G2534,G2535,
G2607,G3330,G2643,G2687,G2725,G2742,G2760,G2794,G2811,G3280,
G3290,G3298,G3316,G3406,G3414,G3422,G1626,G1662,G2567,G2589,
G2608,G2654,G3253,G3277,G3287,G3305,G3313,G3350,G932,G2508,
G2524,G2525,G2526,G3294,G2609,G3410,G3418,G2624,G3426,G2629,
G2647,G2706,G2777,G3264,G3284,G3302,G3303,G3320,G3398,G2657,
G398,G933,G2527,G3259,G3354,G3293,G2563,G3311,G2585,G2625,
G3283,G3286,G3304,G3319,G3322,G3358,G3366,G3382,G3390,G397,
G2544,G2562,G2584,G3402,G2626,G2632,G2634,G2650,G3268,G3256,
G3285,G3321,G3371,G3403,G3411,G362,G1030,G2564,G3362,G3370,
G2586,G3386,G3394,G2633,G3261,G3269,G3347,G3395,G363,G2536,
G3260,G3377,G2580,G3409,G2616,G3417,G2622,G2635,G2805,G2808,
G3334,G3342,G3454,G2537,G3275,G2540,G3353,G2557,G2579,G3401,
G2602,G2615,G2621,G3267,G3112,G3355,G3363,G3379,G3387,G2538,
G2539,G3338,G3346,G2556,G2581,G2601,G2617,G2623,G2638,G3458,
G2814,G2816,G3111,G2541,G2558,G3361,G2571,G3369,G2577,G3385,
G2593,G3393,G2598,G2603,G3113,G3116,G3451,G395,G2570,G2576,
G2592,G2597,G2736,G2739,G2788,G3438,G3446,G3459,G3119,G3120,
G2572,G2578,G2594,G2599,G2677,G3457,G2700,G2771,G3331,G3339,
G3427,G3443,G954,G955,G2600,G3442,G3450,G2676,G2745,G2748,
G3465,G3435,G950,G3337,G2548,G3345,G2553,G2661,G2662,G3433,
G3449,G2672,G2674,G2719,G2754,G3430,G383,G951,G2547,G2552,
G2663,G2670,G3441,G2671,G2675,G3491,G3499,G2549,G2554,G2664,
G3434,G2669,G2673,G2757,G2791,G365,G1031,G2555,G2665,G2667,
G2774,G3497,G3505,G366,G2658,G2659,G2666,G2668,G2681,G2763,
G2765,G2797,G2799,G2660,G2703,G2722,G2780,G2782,G386,G392,
G2684,G3462,G3470,G389,G2709,G2713,G2728,G2730,G2922,G3467,
G2690,G2694,G2821,G3466,G3474,G380,G2822,G3473,G2827,G2839,
G2883,G3507,G2823,G2826,G2880,G2925,G2928,G3510,G2828,G3494,
G3502,G3513,G3544,G3552,G406,G2929,G3475,G3483,G3514,G3515,
G3541,G3549,G2930,G2842,G3498,G2852,G3506,G3548,G3556,G3478,
G3486,G3516,G408,G3481,G3489,G2843,G2853,G3547,G2887,G2896,
G3555,G3520,G2831,G3482,G2836,G3490,G2844,G2848,G2886,G2895,
G2832,G2837,G2849,G3524,G2888,G2891,G2833,G2838,G2892,G3517,
G2906,G2908,G2913,G3523,G2855,G2907,G2909,G3525,G3533,G2854,
G2910,G3560,G3568,G2856,G3539,G3531,G3572,G3564,G3557,G3565,
G3528,G3536,G2921,G2917,G3571,G3563,G2863,G2859,G2920,G2916,
G3540,G3532,G2864,G2860,G403,G404,G400,G401;
buf gate_0(G432,G50);
not gate_1(G442,G50);
buf gate_2(G447,G58);
not gate_3(G456,G58);
buf gate_4(G460,G68);
not gate_5(G463,G68);
buf gate_6(G467,G68);
buf gate_7(G476,G77);
not gate_8(G479,G77);
buf gate_9(G483,G77);
buf gate_10(G492,G87);
not gate_11(G501,G87);
buf gate_12(G504,G97);
not gate_13(G513,G97);
buf gate_14(G517,G107);
not gate_15(G526,G107);
buf gate_16(G530,G116);
not gate_17(G540,G116);
or gate_18(G587,G257,G264);
not gate_19(G704,G1);
buf gate_20(G707,G1);
not gate_21(G714,G1);
buf gate_22(G717,G13);
not gate_23(G724,G13);
and gate_24(G731,G13,G20);
not gate_25(G732,G20);
buf gate_26(G736,G20);
not gate_27(G741,G20);
not gate_28(G758,G33);
buf gate_29(G776,G33);
not gate_30(G780,G33);
and gate_31(G788,G33,G41);
not gate_32(G791,G41);
or gate_33(G798,G41,G45);
buf gate_34(G799,G45);
not gate_35(G802,G45);
not gate_36(G826,G50);
buf gate_37(G828,G58);
not gate_38(G831,G58);
buf gate_39(G833,G68);
not gate_40(G836,G68);
buf gate_41(G839,G87);
not gate_42(G842,G87);
buf gate_43(G845,G97);
not gate_44(G848,G97);
not gate_45(G851,G107);
buf gate_46(G890,G1);
buf gate_47(G898,G68);
buf gate_48(G907,G107);
not gate_49(G1032,G20);
buf gate_50(G1035,G190);
not gate_51(G1048,G200);
and gate_52(G1049,G20,G200);
nand gate_53(G1050,G20,G200);
and gate_54(G1051,G20,G179);
not gate_55(G1540,G20);
or gate_56(G1699,G1698,G33);
nand gate_57(G1826,G1,G13);
nand gate_58(G1827,G1,G20,G33);
not gate_59(G1828,G20);
not gate_60(G2051,G33);
buf gate_61(G2478,G179);
not gate_62(G2865,G213);
buf gate_63(G2868,G343);
buf gate_64(G2931,G226);
buf gate_65(G2934,G232);
buf gate_66(G2939,G238);
buf gate_67(G2942,G244);
buf gate_68(G2947,G250);
buf gate_69(G2950,G257);
buf gate_70(G2957,G264);
buf gate_71(G2960,G270);
buf gate_72(G3007,G50);
buf gate_73(G3079,G58);
buf gate_74(G3087,G58);
buf gate_75(G3095,G97);
buf gate_76(G3103,G97);
buf gate_77(G3419,G330);
and gate_78(G588,G250,G587);
or gate_79(G759,G758,G20);
or gate_80(G1541,G1540,G169);
not gate_81(G1772,G731);
or gate_82(G1829,G1828,G1);
and gate_83(G1834,G1826,G1827);
or gate_84(G2052,G2051,G1);
and gate_85(G625,G826,G831,G836);
nand gate_86(G545,G226,G432);
nand gate_87(G546,G232,G447);
nand gate_88(G547,G238,G467);
nand gate_89(G548,G244,G483);
nand gate_90(G549,G250,G492);
nand gate_91(G550,G257,G504);
nand gate_92(G551,G264,G517);
nand gate_93(G552,G270,G530);
not gate_94(G2937,G2931);
not gate_95(G2938,G2934);
not gate_96(G2945,G2939);
not gate_97(G2946,G2942);
nand gate_98(G621,G456,G463);
nand gate_99(G626,G513,G526);
nand gate_100(G635,G460,G476);
buf gate_101(G636,G442);
not gate_102(G3085,G3079);
not gate_103(G3101,G3095);
buf gate_104(G657,G802);
buf gate_105(G675,G802);
buf gate_106(G721,G717);
buf gate_107(G784,G780);
buf gate_108(G794,G791);
and gate_109(G807,G714,G798);
and gate_110(G816,G714,G799,G791);
and gate_111(G823,G704,G799);
and gate_112(G860,G707,G724,G736);
nand gate_113(G861,G707,G724,G736);
nand gate_114(G864,G707,G724);
buf gate_115(G893,G890);
nand gate_116(G896,G717,G732,G45);
nand gate_117(G897,G826,G831,G836);
not gate_118(G3093,G3087);
and gate_119(G905,G842,G848,G851);
nand gate_120(G906,G842,G848,G851);
not gate_121(G3109,G3103);
not gate_122(G973,G741);
not gate_123(G980,G741);
not gate_124(G987,G741);
not gate_125(G994,G741);
not gate_126(G1001,G741);
not gate_127(G1008,G741);
not gate_128(G1015,G741);
not gate_129(G1022,G741);
or gate_130(G1038,G1032,G1035);
nor gate_131(G1043,G1032,G1035);
buf gate_132(G1054,G1051);
not gate_133(G1057,G1051);
buf gate_134(G1512,G776);
buf gate_135(G1681,G780);
not gate_136(G1717,G1699);
not gate_137(G1724,G1699);
not gate_138(G1731,G1699);
not gate_139(G1738,G1699);
not gate_140(G1745,G1699);
not gate_141(G1752,G1699);
not gate_142(G1759,G1699);
not gate_143(G1766,G1699);
or gate_144(G1773,G1,G1772);
not gate_145(G1790,G788);
not gate_146(G1808,G788);
and gate_147(G2278,G704,G717,G732);
not gate_148(G2481,G2478);
not gate_149(G3425,G3419);
or gate_150(G2871,G2865,G2868);
nor gate_151(G2874,G2865,G2868);
not gate_152(G2953,G2947);
not gate_153(G2954,G2950);
not gate_154(G2963,G2957);
not gate_155(G2964,G2960);
buf gate_156(G3010,G456);
not gate_157(G3013,G3007);
buf gate_158(G3017,G463);
buf gate_159(G3020,G479);
buf gate_160(G3027,G501);
buf gate_161(G3030,G513);
buf gate_162(G3037,G526);
buf gate_163(G3040,G540);
buf gate_164(G3082,G898);
buf gate_165(G3090,G898);
buf gate_166(G3098,G907);
buf gate_167(G3106,G907);
nand gate_168(G352,G479,G625);
and gate_169(G553,G545,G546,G547,G548);
and gate_170(G554,G549,G550,G551,G552);
nand gate_171(G555,G2934,G2937);
nand gate_172(G556,G2931,G2938);
nand gate_173(G560,G2942,G2945);
nand gate_174(G561,G2939,G2946);
and gate_175(G650,G432,G621);
and gate_176(G956,G890,G896);
not gate_177(G974,G759);
and gate_178(G975,G741,G759);
and gate_179(G976,G897,G973);
not gate_180(G981,G759);
and gate_181(G982,G741,G759);
not gate_182(G988,G759);
and gate_183(G989,G741,G759);
and gate_184(G990,G836,G987);
not gate_185(G995,G759);
and gate_186(G996,G741,G759);
and gate_187(G997,G77,G994);
not gate_188(G1002,G759);
and gate_189(G1003,G741,G759);
and gate_190(G1004,G906,G1001);
not gate_191(G1009,G759);
and gate_192(G1010,G741,G759);
not gate_193(G1016,G759);
and gate_194(G1017,G741,G759);
and gate_195(G1018,G851,G1015);
not gate_196(G1023,G759);
and gate_197(G1024,G741,G759);
and gate_198(G1025,G116,G1022);
and gate_199(G1720,G222,G1717);
and gate_200(G1727,G223,G1724);
and gate_201(G1734,G226,G1731);
and gate_202(G1741,G232,G1738);
and gate_203(G1748,G238,G1745);
and gate_204(G1755,G244,G1752);
and gate_205(G1762,G250,G1759);
and gate_206(G1769,G257,G1766);
and gate_207(G1791,G1,G13,G1790);
and gate_208(G1809,G1,G13,G1808);
not gate_209(G1851,G1834);
not gate_210(G1901,G1834);
not gate_211(G1952,G1834);
not gate_212(G2002,G1834);
not gate_213(G2057,G1834);
not gate_214(G2109,G1834);
not gate_215(G2162,G1834);
not gate_216(G2214,G1834);
nand gate_217(G2955,G2950,G2953);
nand gate_218(G2956,G2947,G2954);
nand gate_219(G2965,G2960,G2963);
nand gate_220(G2966,G2957,G2964);
not gate_221(G353,G352);
and gate_222(G354,G87,G626);
nand gate_223(G557,G555,G556);
nand gate_224(G562,G560,G561);
nand gate_225(G586,G553,G554);
and gate_226(G630,G540,G905);
nand gate_227(G634,G540,G905);
not gate_228(G639,G636);
nand gate_229(G642,G3082,G3085);
not gate_230(G3086,G3082);
and gate_231(G644,G460,G636);
nand gate_232(G646,G3098,G3101);
not gate_233(G3102,G3098);
nand gate_234(G654,G87,G626);
not gate_235(G660,G657);
not gate_236(G678,G675);
nand gate_237(G804,G860,G776);
nand gate_238(G806,G860,G780);
nand gate_239(G855,G707,G721,G736);
nand gate_240(G867,G707,G724,G736,G794);
nand gate_241(G903,G3090,G3093);
not gate_242(G3094,G3090);
nand gate_243(G912,G3106,G3109);
not gate_244(G3110,G3106);
not gate_245(G915,G861);
not gate_246(G927,G893);
not gate_247(G941,G864);
and gate_248(G977,G828,G974);
and gate_249(G978,G150,G975);
and gate_250(G984,G833,G981);
and gate_251(G985,G159,G982);
and gate_252(G991,G77,G988);
and gate_253(G992,G50,G989);
and gate_254(G998,G839,G995);
and gate_255(G999,G828,G996);
and gate_256(G1005,G845,G1002);
and gate_257(G1006,G833,G1003);
and gate_258(G1012,G107,G1009);
and gate_259(G1013,G77,G1010);
and gate_260(G1019,G116,G1016);
and gate_261(G1020,G839,G1017);
and gate_262(G1026,G283,G1023);
and gate_263(G1027,G845,G1024);
and gate_264(G1060,G200,G1054);
and gate_265(G1063,G1048,G1054);
and gate_266(G1066,G1049,G1057);
and gate_267(G1069,G1050,G1057);
nand gate_268(G1527,G784,G794);
nand gate_269(G1530,G776,G794);
nand gate_270(G1542,G707,G721,G1541);
nand gate_271(G1563,G724,G732,G784);
nand gate_272(G1572,G724,G784);
not gate_273(G1581,G1512);
not gate_274(G1585,G1512);
not gate_275(G1589,G1512);
not gate_276(G1593,G1512);
not gate_277(G1597,G1512);
not gate_278(G1601,G1512);
not gate_279(G1605,G1512);
not gate_280(G1716,G1681);
and gate_281(G1718,G1681,G1699);
not gate_282(G1723,G1681);
and gate_283(G1725,G1681,G1699);
not gate_284(G1730,G1681);
and gate_285(G1732,G1681,G1699);
not gate_286(G1737,G1681);
and gate_287(G1739,G1681,G1699);
not gate_288(G1744,G1681);
and gate_289(G1746,G1681,G1699);
not gate_290(G1751,G1681);
and gate_291(G1753,G1681,G1699);
not gate_292(G1758,G1681);
and gate_293(G1760,G1681,G1699);
not gate_294(G1765,G1681);
and gate_295(G1767,G1681,G1699);
and gate_296(G1852,G1834,G1773);
nor gate_297(G1856,G50,G1773);
not gate_298(G1870,G807);
and gate_299(G1902,G1834,G1773);
nor gate_300(G1906,G58,G1773);
not gate_301(G1920,G807);
and gate_302(G1953,G1834,G1773);
nor gate_303(G1957,G68,G1773);
not gate_304(G1971,G807);
and gate_305(G2003,G1834,G1773);
nor gate_306(G2007,G77,G1773);
not gate_307(G2021,G807);
and gate_308(G2058,G1834,G1773);
nor gate_309(G2062,G87,G1773);
not gate_310(G2076,G823);
and gate_311(G2110,G1834,G1773);
nor gate_312(G2114,G97,G1773);
not gate_313(G2128,G816);
and gate_314(G2163,G1834,G1773);
nor gate_315(G2167,G107,G1773);
not gate_316(G2181,G816);
and gate_317(G2215,G1834,G1773);
nor gate_318(G2219,G116,G1773);
not gate_319(G2233,G816);
and gate_320(G2285,G2278,G213);
nand gate_321(G2288,G2278,G213);
and gate_322(G2289,G2278,G213,G343);
nand gate_323(G2293,G2278,G213,G343);
and gate_324(G2298,G2278,G213,G343);
nand gate_325(G2302,G2278,G213,G343);
buf gate_326(G2877,G2874);
nand gate_327(G2983,G2955,G2956);
nand gate_328(G2986,G2965,G2966);
not gate_329(G3014,G3010);
nand gate_330(G3015,G3010,G3013);
not gate_331(G3023,G3017);
not gate_332(G3024,G3020);
not gate_333(G3033,G3027);
not gate_334(G3034,G3030);
not gate_335(G3043,G3037);
not gate_336(G3044,G3040);
not gate_337(G355,G354);
nand gate_338(G643,G3079,G3086);
nand gate_339(G647,G3095,G3102);
and gate_340(G680,G650,G675);
nand gate_341(G904,G3087,G3094);
nand gate_342(G913,G3103,G3110);
and gate_343(G920,G588,G915);
or gate_344(G979,G976,G977,G978);
or gate_345(G993,G990,G991,G992);
or gate_346(G1000,G997,G998,G999);
or gate_347(G1007,G1004,G1005,G1006);
or gate_348(G1021,G1018,G1019,G1020);
or gate_349(G1028,G1025,G1026,G1027);
and gate_350(G1719,G77,G1716);
and gate_351(G1721,G223,G1718);
and gate_352(G1726,G87,G1723);
and gate_353(G1728,G226,G1725);
and gate_354(G1733,G97,G1730);
and gate_355(G1735,G232,G1732);
and gate_356(G1740,G107,G1737);
and gate_357(G1742,G238,G1739);
and gate_358(G1747,G116,G1744);
and gate_359(G1749,G244,G1746);
and gate_360(G1754,G283,G1751);
and gate_361(G1756,G250,G1753);
and gate_362(G1761,G294,G1758);
and gate_363(G1763,G257,G1760);
and gate_364(G1768,G303,G1765);
and gate_365(G1770,G264,G1767);
buf gate_366(G1794,G1791);
not gate_367(G1799,G1791);
buf gate_368(G1812,G1809);
not gate_369(G1817,G1809);
and gate_370(G1859,G50,G1829,G1852);
and gate_371(G1909,G58,G1829,G1902);
and gate_372(G1960,G68,G1829,G1953);
and gate_373(G2010,G77,G1829,G2003);
and gate_374(G2065,G87,G2052,G2058);
and gate_375(G2117,G97,G2052,G2110);
and gate_376(G2170,G107,G2052,G2163);
and gate_377(G2222,G116,G2052,G2215);
not gate_378(G2678,G956);
not gate_379(G2697,G956);
not gate_380(G2716,G956);
not gate_381(G2733,G956);
not gate_382(G2751,G956);
not gate_383(G2768,G956);
not gate_384(G2785,G956);
not gate_385(G2802,G956);
nand gate_386(G3016,G3007,G3014);
nand gate_387(G3025,G3020,G3023);
nand gate_388(G3026,G3017,G3024);
nand gate_389(G3035,G3030,G3033);
nand gate_390(G3036,G3027,G3034);
nand gate_391(G3045,G3040,G3043);
nand gate_392(G3046,G3037,G3044);
not gate_393(G2989,G2983);
not gate_394(G2990,G2986);
not gate_395(G610,G804);
and gate_396(G613,G804,G806);
not gate_397(G616,G806);
nand gate_398(G640,G642,G643);
nand gate_399(G648,G646,G647);
and gate_400(G655,G630,G635,G442,G58);
not gate_401(G665,G804);
and gate_402(G668,G804,G806);
not gate_403(G671,G806);
not gate_404(G683,G804);
not gate_405(G685,G806);
and gate_406(G688,G804,G806);
not gate_407(G694,G804);
not gate_408(G696,G806);
and gate_409(G699,G804,G806);
buf gate_410(G870,G867);
buf gate_411(G887,G867);
nand gate_412(G901,G903,G904);
nand gate_413(G910,G912,G913);
not gate_414(G914,G855);
and gate_415(G916,G855,G861);
not gate_416(G942,G855);
and gate_417(G943,G864,G855);
nand gate_418(G1072,G1043,G1069);
nand gate_419(G1084,G1043,G1066);
nand gate_420(G1096,G1038,G1069);
nand gate_421(G1108,G1038,G1066);
nand gate_422(G1120,G1043,G1063);
nand gate_423(G1132,G1043,G1060);
nand gate_424(G1144,G1038,G1063);
nand gate_425(G1156,G1038,G1060);
not gate_426(G1533,G1527);
not gate_427(G1534,G1530);
and gate_428(G1535,G1527,G1530);
buf gate_429(G1545,G1542);
buf gate_430(G1554,G1542);
not gate_431(G1610,G1572);
not gate_432(G1619,G1572);
not gate_433(G1628,G1572);
not gate_434(G1637,G1572);
not gate_435(G1646,G1563);
not gate_436(G1655,G1563);
not gate_437(G1664,G1563);
not gate_438(G1673,G1563);
or gate_439(G1722,G1719,G1720,G1721);
or gate_440(G1729,G1726,G1727,G1728);
or gate_441(G1736,G1733,G1734,G1735);
or gate_442(G1743,G1740,G1741,G1742);
or gate_443(G1750,G1747,G1748,G1749);
or gate_444(G1757,G1754,G1755,G1756);
or gate_445(G1764,G1761,G1762,G1763);
or gate_446(G1771,G1768,G1769,G1770);
and gate_447(G1853,G979,G1851);
and gate_448(G1954,G993,G1952);
and gate_449(G2004,G1000,G2002);
and gate_450(G2059,G1007,G2057);
and gate_451(G2164,G1021,G2162);
and gate_452(G2216,G1028,G2214);
buf gate_453(G2485,G2293);
and gate_454(G2900,G2877,G2897);
nand gate_455(G2903,G2877,G2897);
buf gate_456(G2967,G557);
buf gate_457(G2970,G562);
buf gate_458(G2975,G557);
buf gate_459(G2978,G562);
nand gate_460(G3047,G3015,G3016);
nand gate_461(G3050,G3025,G3026);
nand gate_462(G3055,G3035,G3036);
nand gate_463(G3058,G3045,G3046);
nand gate_464(G574,G2986,G2989);
nand gate_465(G575,G2983,G2990);
and gate_466(G617,G501,G613);
and gate_467(G641,G640,G476,G639);
and gate_468(G649,G530,G648);
and gate_469(G662,G655,G657);
and gate_470(G672,G513,G668);
and gate_471(G690,G654,G685);
and gate_472(G691,G540,G688);
and gate_473(G701,G634,G696);
and gate_474(G702,G526,G699);
not gate_475(G902,G901);
not gate_476(G911,G910);
and gate_477(G917,G650,G914);
and gate_478(G923,G586,G916);
and gate_479(G1538,G442,G1535);
and gate_480(G1871,G1817,G226,G1870);
and gate_481(G1872,G1817,G274,G807);
and gate_482(G1873,G1812,G1722);
and gate_483(G1921,G1817,G232,G1920);
and gate_484(G1922,G1817,G274,G807);
and gate_485(G1923,G1812,G1729);
and gate_486(G1972,G1817,G238,G1971);
and gate_487(G1973,G1817,G274,G807);
and gate_488(G1974,G1812,G1736);
and gate_489(G2022,G1817,G244,G2021);
and gate_490(G2023,G1817,G274,G807);
and gate_491(G2024,G1812,G1743);
and gate_492(G2077,G1799,G250,G2076);
and gate_493(G2078,G1799,G274,G823);
and gate_494(G2079,G1794,G1750);
and gate_495(G2129,G1799,G257,G2128);
and gate_496(G2130,G1799,G274,G816);
and gate_497(G2131,G1794,G1757);
and gate_498(G2182,G1799,G264,G2181);
and gate_499(G2183,G1799,G274,G816);
and gate_500(G2184,G1794,G1764);
and gate_501(G2234,G1799,G270,G2233);
and gate_502(G2235,G1799,G274,G816);
and gate_503(G2236,G1794,G1771);
not gate_504(G2973,G2967);
not gate_505(G2974,G2970);
not gate_506(G2981,G2975);
not gate_507(G2982,G2978);
nand gate_508(G576,G574,G575);
not gate_509(G3053,G3047);
not gate_510(G3054,G3050);
not gate_511(G3061,G3055);
not gate_512(G3062,G3058);
or gate_513(G645,G641,G644);
not gate_514(G926,G887);
and gate_515(G928,G887,G893);
and gate_516(G947,G649,G942);
and gate_517(G983,G902,G980);
and gate_518(G1011,G911,G1008);
buf gate_519(G1075,G1072);
buf gate_520(G1087,G1084);
buf gate_521(G1099,G1096);
buf gate_522(G1111,G1108);
buf gate_523(G1123,G1120);
buf gate_524(G1135,G1132);
buf gate_525(G1147,G1144);
buf gate_526(G1159,G1156);
buf gate_527(G1168,G1072);
buf gate_528(G1177,G1084);
buf gate_529(G1186,G1096);
buf gate_530(G1195,G1108);
buf gate_531(G1204,G1120);
buf gate_532(G1213,G1132);
buf gate_533(G1222,G1144);
buf gate_534(G1231,G1156);
not gate_535(G1609,G1545);
and gate_536(G1611,G1545,G1572);
not gate_537(G1618,G1545);
and gate_538(G1620,G1545,G1572);
not gate_539(G1627,G1545);
and gate_540(G1629,G1545,G1572);
not gate_541(G1636,G1545);
and gate_542(G1638,G1545,G1572);
not gate_543(G1645,G1554);
and gate_544(G1647,G1554,G1563);
not gate_545(G1654,G1554);
and gate_546(G1656,G1554,G1563);
not gate_547(G1663,G1554);
and gate_548(G1665,G1554,G1563);
not gate_549(G1672,G1554);
and gate_550(G1674,G1554,G1563);
or gate_551(G1862,G1853,G1856,G1859);
nor gate_552(G1866,G1853,G1856,G1859);
or gate_553(G1874,G1871,G1872,G1873);
or gate_554(G1924,G1921,G1922,G1923);
or gate_555(G1963,G1954,G1957,G1960);
nor gate_556(G1967,G1954,G1957,G1960);
or gate_557(G1975,G1972,G1973,G1974);
or gate_558(G2013,G2004,G2007,G2010);
nor gate_559(G2017,G2004,G2007,G2010);
or gate_560(G2025,G2022,G2023,G2024);
or gate_561(G2068,G2059,G2062,G2065);
nor gate_562(G2072,G2059,G2062,G2065);
or gate_563(G2080,G2077,G2078,G2079);
or gate_564(G2132,G2129,G2130,G2131);
or gate_565(G2173,G2164,G2167,G2170);
nor gate_566(G2177,G2164,G2167,G2170);
or gate_567(G2185,G2182,G2183,G2184);
or gate_568(G2225,G2216,G2219,G2222);
nor gate_569(G2229,G2216,G2219,G2222);
or gate_570(G2237,G2234,G2235,G2236);
not gate_571(G2488,G2485);
not gate_572(G2679,G870);
and gate_573(G2680,G956,G870);
not gate_574(G2698,G870);
and gate_575(G2699,G956,G870);
not gate_576(G2717,G870);
and gate_577(G2718,G956,G870);
not gate_578(G2734,G870);
and gate_579(G2735,G956,G870);
not gate_580(G2752,G870);
and gate_581(G2753,G956,G870);
not gate_582(G2769,G870);
and gate_583(G2770,G956,G870);
not gate_584(G2786,G870);
and gate_585(G2787,G956,G870);
not gate_586(G2803,G870);
and gate_587(G2804,G956,G870);
or gate_588(G359,G917,G920,G923);
nor gate_589(G1029,G917,G920,G923);
nand gate_590(G565,G2970,G2973);
nand gate_591(G566,G2967,G2974);
nand gate_592(G569,G2978,G2981);
nand gate_593(G570,G2975,G2982);
nand gate_594(G589,G3050,G3053);
nand gate_595(G590,G3047,G3054);
nand gate_596(G595,G3058,G3061);
nand gate_597(G596,G3055,G3062);
and gate_598(G929,G650,G926);
and gate_599(G938,G630,G928);
and gate_600(G944,G645,G941);
or gate_601(G986,G983,G984,G985);
or gate_602(G1014,G1011,G1012,G1013);
and gate_603(G1616,G442,G1611);
and gate_604(G1625,G456,G1620);
and gate_605(G1634,G463,G1629);
and gate_606(G1643,G479,G1638);
not gate_607(G360,G1029);
nand gate_608(G567,G565,G566);
nand gate_609(G571,G569,G570);
buf gate_610(G579,G576);
nand gate_611(G591,G589,G590);
nand gate_612(G597,G595,G596);
and gate_613(G614,G576,G610);
not gate_614(G1240,G1075);
not gate_615(G1241,G1087);
not gate_616(G1242,G1099);
not gate_617(G1243,G1111);
not gate_618(G1244,G1123);
not gate_619(G1245,G1135);
not gate_620(G1246,G1147);
not gate_621(G1247,G1159);
not gate_622(G1257,G1075);
not gate_623(G1258,G1087);
not gate_624(G1259,G1099);
not gate_625(G1260,G1111);
not gate_626(G1261,G1123);
not gate_627(G1262,G1135);
not gate_628(G1263,G1147);
not gate_629(G1264,G1159);
not gate_630(G1274,G1075);
not gate_631(G1275,G1087);
not gate_632(G1276,G1099);
not gate_633(G1277,G1111);
not gate_634(G1278,G1123);
not gate_635(G1279,G1135);
not gate_636(G1280,G1147);
not gate_637(G1281,G1159);
not gate_638(G1291,G1075);
not gate_639(G1292,G1087);
not gate_640(G1293,G1099);
not gate_641(G1294,G1111);
not gate_642(G1295,G1123);
not gate_643(G1296,G1135);
not gate_644(G1297,G1147);
not gate_645(G1298,G1159);
not gate_646(G1308,G1075);
not gate_647(G1309,G1087);
not gate_648(G1310,G1099);
not gate_649(G1311,G1111);
not gate_650(G1312,G1123);
not gate_651(G1313,G1135);
not gate_652(G1314,G1147);
not gate_653(G1315,G1159);
not gate_654(G1325,G1075);
not gate_655(G1326,G1087);
not gate_656(G1327,G1099);
not gate_657(G1328,G1111);
not gate_658(G1329,G1123);
not gate_659(G1330,G1135);
not gate_660(G1331,G1147);
not gate_661(G1332,G1159);
not gate_662(G1342,G1075);
not gate_663(G1343,G1087);
not gate_664(G1344,G1099);
not gate_665(G1345,G1111);
not gate_666(G1346,G1123);
not gate_667(G1347,G1135);
not gate_668(G1348,G1147);
not gate_669(G1349,G1159);
not gate_670(G1359,G1075);
not gate_671(G1360,G1087);
not gate_672(G1361,G1099);
not gate_673(G1362,G1111);
not gate_674(G1363,G1123);
not gate_675(G1364,G1135);
not gate_676(G1365,G1147);
not gate_677(G1366,G1159);
not gate_678(G1376,G1168);
not gate_679(G1377,G1177);
not gate_680(G1378,G1186);
not gate_681(G1379,G1195);
not gate_682(G1380,G1204);
not gate_683(G1381,G1213);
not gate_684(G1382,G1222);
not gate_685(G1383,G1231);
not gate_686(G1393,G1168);
not gate_687(G1394,G1177);
not gate_688(G1395,G1186);
not gate_689(G1396,G1195);
not gate_690(G1397,G1204);
not gate_691(G1398,G1213);
not gate_692(G1399,G1222);
not gate_693(G1400,G1231);
not gate_694(G1410,G1168);
not gate_695(G1411,G1177);
not gate_696(G1412,G1186);
not gate_697(G1413,G1195);
not gate_698(G1414,G1204);
not gate_699(G1415,G1213);
not gate_700(G1416,G1222);
not gate_701(G1417,G1231);
not gate_702(G1427,G1168);
not gate_703(G1428,G1177);
not gate_704(G1429,G1186);
not gate_705(G1430,G1195);
not gate_706(G1431,G1204);
not gate_707(G1432,G1213);
not gate_708(G1433,G1222);
not gate_709(G1434,G1231);
not gate_710(G1444,G1168);
not gate_711(G1445,G1177);
not gate_712(G1446,G1186);
not gate_713(G1447,G1195);
not gate_714(G1448,G1204);
not gate_715(G1449,G1213);
not gate_716(G1450,G1222);
not gate_717(G1451,G1231);
not gate_718(G1461,G1168);
not gate_719(G1462,G1177);
not gate_720(G1463,G1186);
not gate_721(G1464,G1195);
not gate_722(G1465,G1204);
not gate_723(G1466,G1213);
not gate_724(G1467,G1222);
not gate_725(G1468,G1231);
not gate_726(G1478,G1168);
not gate_727(G1479,G1177);
not gate_728(G1480,G1186);
not gate_729(G1481,G1195);
not gate_730(G1482,G1204);
not gate_731(G1483,G1213);
not gate_732(G1484,G1222);
not gate_733(G1485,G1231);
not gate_734(G1495,G1168);
not gate_735(G1496,G1177);
not gate_736(G1497,G1186);
not gate_737(G1498,G1195);
not gate_738(G1499,G1204);
not gate_739(G1500,G1213);
not gate_740(G1501,G1222);
not gate_741(G1502,G1231);
buf gate_742(G1877,G1874);
not gate_743(G1880,G1874);
not gate_744(G1891,G1866);
and gate_745(G1903,G986,G1901);
buf gate_746(G1927,G1924);
not gate_747(G1930,G1924);
buf gate_748(G1978,G1975);
not gate_749(G1981,G1975);
not gate_750(G1992,G1967);
buf gate_751(G2028,G2025);
not gate_752(G2031,G2025);
not gate_753(G2042,G2017);
buf gate_754(G2085,G2080);
not gate_755(G2088,G2080);
not gate_756(G2099,G2072);
and gate_757(G2111,G1014,G2109);
buf gate_758(G2137,G2132);
not gate_759(G2140,G2132);
buf gate_760(G2190,G2185);
not gate_761(G2193,G2185);
not gate_762(G2204,G2177);
buf gate_763(G2242,G2237);
not gate_764(G2245,G2237);
not gate_765(G2256,G2229);
and gate_766(G2320,G2285,G1862);
and gate_767(G2341,G2289,G1963);
and gate_768(G2354,G2289,G2013);
and gate_769(G2367,G2289,G2068);
and gate_770(G2383,G2298,G2173);
and gate_771(G2391,G2298,G2225);
not gate_772(G2474,G2080);
not gate_773(G2475,G2132);
not gate_774(G2476,G2185);
not gate_775(G2477,G2237);
and gate_776(G2482,G2080,G2132,G2185,G2237,G2481);
nand gate_777(G361,G359,G360);
not gate_778(G568,G567);
or gate_779(G618,G614,G616,G617);
and gate_780(G1248,G124,G1240);
and gate_781(G1249,G159,G1241);
and gate_782(G1250,G150,G1242);
and gate_783(G1251,G143,G1243);
and gate_784(G1252,G137,G1244);
and gate_785(G1253,G132,G1245);
and gate_786(G1254,G128,G1246);
and gate_787(G1255,G125,G1247);
and gate_788(G1265,G125,G1257);
and gate_789(G1266,G432,G1258);
and gate_790(G1267,G159,G1259);
and gate_791(G1268,G150,G1260);
and gate_792(G1269,G143,G1261);
and gate_793(G1270,G137,G1262);
and gate_794(G1271,G132,G1263);
and gate_795(G1272,G128,G1264);
and gate_796(G1282,G128,G1274);
and gate_797(G1283,G447,G1275);
and gate_798(G1284,G432,G1276);
and gate_799(G1285,G159,G1277);
and gate_800(G1286,G150,G1278);
and gate_801(G1287,G143,G1279);
and gate_802(G1288,G137,G1280);
and gate_803(G1289,G132,G1281);
and gate_804(G1299,G132,G1291);
and gate_805(G1300,G467,G1292);
and gate_806(G1301,G447,G1293);
and gate_807(G1302,G432,G1294);
and gate_808(G1303,G159,G1295);
and gate_809(G1304,G150,G1296);
and gate_810(G1305,G143,G1297);
and gate_811(G1306,G137,G1298);
and gate_812(G1316,G137,G1308);
and gate_813(G1317,G483,G1309);
and gate_814(G1318,G467,G1310);
and gate_815(G1319,G447,G1311);
and gate_816(G1320,G432,G1312);
and gate_817(G1321,G159,G1313);
and gate_818(G1322,G150,G1314);
and gate_819(G1323,G143,G1315);
and gate_820(G1333,G143,G1325);
and gate_821(G1334,G492,G1326);
and gate_822(G1335,G483,G1327);
and gate_823(G1336,G467,G1328);
and gate_824(G1337,G447,G1329);
and gate_825(G1338,G432,G1330);
and gate_826(G1339,G159,G1331);
and gate_827(G1340,G150,G1332);
and gate_828(G1350,G150,G1342);
and gate_829(G1351,G504,G1343);
and gate_830(G1352,G492,G1344);
and gate_831(G1353,G483,G1345);
and gate_832(G1354,G467,G1346);
and gate_833(G1355,G447,G1347);
and gate_834(G1356,G432,G1348);
and gate_835(G1357,G159,G1349);
and gate_836(G1367,G159,G1359);
and gate_837(G1368,G517,G1360);
and gate_838(G1369,G504,G1361);
and gate_839(G1370,G492,G1362);
and gate_840(G1371,G483,G1363);
and gate_841(G1372,G467,G1364);
and gate_842(G1373,G447,G1365);
and gate_843(G1374,G432,G1366);
and gate_844(G1384,G283,G1376);
and gate_845(G1385,G447,G1377);
and gate_846(G1386,G467,G1378);
and gate_847(G1387,G483,G1379);
and gate_848(G1388,G492,G1380);
and gate_849(G1389,G504,G1381);
and gate_850(G1390,G517,G1382);
and gate_851(G1391,G530,G1383);
and gate_852(G1401,G294,G1393);
and gate_853(G1402,G467,G1394);
and gate_854(G1403,G483,G1395);
and gate_855(G1404,G492,G1396);
and gate_856(G1405,G504,G1397);
and gate_857(G1406,G517,G1398);
and gate_858(G1407,G530,G1399);
and gate_859(G1408,G283,G1400);
and gate_860(G1418,G303,G1410);
and gate_861(G1419,G483,G1411);
and gate_862(G1420,G492,G1412);
and gate_863(G1421,G504,G1413);
and gate_864(G1422,G517,G1414);
and gate_865(G1423,G530,G1415);
and gate_866(G1424,G283,G1416);
and gate_867(G1425,G294,G1417);
and gate_868(G1435,G311,G1427);
and gate_869(G1436,G492,G1428);
and gate_870(G1437,G504,G1429);
and gate_871(G1438,G517,G1430);
and gate_872(G1439,G530,G1431);
and gate_873(G1440,G283,G1432);
and gate_874(G1441,G294,G1433);
and gate_875(G1442,G303,G1434);
and gate_876(G1452,G317,G1444);
and gate_877(G1453,G504,G1445);
and gate_878(G1454,G517,G1446);
and gate_879(G1455,G530,G1447);
and gate_880(G1456,G283,G1448);
and gate_881(G1457,G294,G1449);
and gate_882(G1458,G303,G1450);
and gate_883(G1459,G311,G1451);
and gate_884(G1469,G322,G1461);
and gate_885(G1470,G517,G1462);
and gate_886(G1471,G530,G1463);
and gate_887(G1472,G283,G1464);
and gate_888(G1473,G294,G1465);
and gate_889(G1474,G303,G1466);
and gate_890(G1475,G311,G1467);
and gate_891(G1476,G317,G1468);
and gate_892(G1486,G326,G1478);
and gate_893(G1487,G530,G1479);
and gate_894(G1488,G283,G1480);
and gate_895(G1489,G294,G1481);
and gate_896(G1490,G303,G1482);
and gate_897(G1491,G311,G1483);
and gate_898(G1492,G317,G1484);
and gate_899(G1493,G322,G1485);
and gate_900(G1503,G329,G1495);
and gate_901(G1504,G283,G1496);
and gate_902(G1505,G294,G1497);
and gate_903(G1506,G303,G1498);
and gate_904(G1507,G311,G1499);
and gate_905(G1508,G317,G1500);
and gate_906(G1509,G322,G1501);
and gate_907(G1510,G326,G1502);
and gate_908(G2483,G2474,G2475,G2476,G2477,G2478);
buf gate_909(G600,G597);
and gate_910(G661,G568,G660);
and gate_911(G669,G597,G665);
and gate_912(G679,G591,G678);
nor gate_913(G1256,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255);
nor gate_914(G1273,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272);
nor gate_915(G1290,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289);
nor gate_916(G1307,G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306);
nor gate_917(G1324,G1316,G1317,G1318,G1319,G1320,G1321,G1322,G1323);
nor gate_918(G1341,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340);
nor gate_919(G1358,G1350,G1351,G1352,G1353,G1354,G1355,G1356,G1357);
nor gate_920(G1375,G1367,G1368,G1369,G1370,G1371,G1372,G1373,G1374);
nor gate_921(G1392,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391);
nor gate_922(G1409,G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408);
nor gate_923(G1426,G1418,G1419,G1420,G1421,G1422,G1423,G1424,G1425);
nor gate_924(G1443,G1435,G1436,G1437,G1438,G1439,G1440,G1441,G1442);
nor gate_925(G1460,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459);
nor gate_926(G1477,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476);
nor gate_927(G1494,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493);
nor gate_928(G1511,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510);
and gate_929(G1652,G618,G1647);
and gate_930(G1883,G169,G1862,G1877);
and gate_931(G1886,G179,G1862,G1880);
and gate_932(G1889,G190,G1866,G1880);
and gate_933(G1890,G200,G1866,G1877);
or gate_934(G1912,G1903,G1906,G1909);
nor gate_935(G1916,G1903,G1906,G1909);
and gate_936(G1984,G169,G1963,G1978);
and gate_937(G1987,G179,G1963,G1981);
and gate_938(G1990,G190,G1967,G1981);
and gate_939(G1991,G200,G1967,G1978);
and gate_940(G2034,G169,G2013,G2028);
and gate_941(G2037,G179,G2013,G2031);
and gate_942(G2040,G190,G2017,G2031);
and gate_943(G2041,G200,G2017,G2028);
and gate_944(G2091,G169,G2068,G2085);
and gate_945(G2094,G179,G2068,G2088);
and gate_946(G2097,G190,G2072,G2088);
and gate_947(G2098,G200,G2072,G2085);
or gate_948(G2120,G2111,G2114,G2117);
nor gate_949(G2124,G2111,G2114,G2117);
and gate_950(G2196,G169,G2173,G2190);
and gate_951(G2199,G179,G2173,G2193);
and gate_952(G2202,G190,G2177,G2193);
and gate_953(G2203,G200,G2177,G2190);
and gate_954(G2248,G169,G2225,G2242);
and gate_955(G2251,G179,G2225,G2245);
and gate_956(G2254,G190,G2229,G2245);
and gate_957(G2255,G200,G2229,G2242);
or gate_958(G2484,G2482,G2483);
buf gate_959(G2991,G571);
buf gate_960(G2994,G579);
buf gate_961(G2999,G571);
buf gate_962(G3002,G579);
buf gate_963(G3063,G591);
buf gate_964(G3071,G591);
buf gate_965(G3124,G2320);
buf gate_966(G3134,G2320);
buf gate_967(G3158,G2341);
buf gate_968(G3166,G2341);
buf gate_969(G3174,G2354);
buf gate_970(G3182,G2354);
buf gate_971(G3190,G2367);
buf gate_972(G3200,G2367);
buf gate_973(G3224,G2383);
buf gate_974(G3232,G2383);
buf gate_975(G3240,G2391);
buf gate_976(G3248,G2391);
nor gate_977(G663,G661,G662);
or gate_978(G673,G669,G671,G672);
nor gate_979(G681,G679,G680);
and gate_980(G1536,G1256,G1533);
and gate_981(G1537,G1392,G1534);
and gate_982(G1582,G1273,G1581);
and gate_983(G1583,G1409,G1512);
and gate_984(G1586,G1290,G1585);
and gate_985(G1587,G1426,G1512);
and gate_986(G1590,G1307,G1589);
and gate_987(G1591,G1443,G1512);
and gate_988(G1594,G1324,G1593);
and gate_989(G1595,G1460,G1512);
and gate_990(G1598,G1341,G1597);
and gate_991(G1599,G1477,G1512);
and gate_992(G1602,G1358,G1601);
and gate_993(G1603,G1494,G1512);
and gate_994(G1606,G1375,G1605);
and gate_995(G1607,G1511,G1512);
or gate_996(G1894,G1889,G1890,G1891);
or gate_997(G1997,G1990,G1991,G1992);
or gate_998(G2047,G2040,G2041,G2042);
or gate_999(G2102,G2097,G2098,G2099);
or gate_1000(G2209,G2202,G2203,G2204);
or gate_1001(G2261,G2254,G2255,G2256);
and gate_1002(G2489,G2484,G2488);
not gate_1003(G3005,G2999);
not gate_1004(G3006,G3002);
not gate_1005(G3077,G3071);
not gate_1006(G3069,G3063);
not gate_1007(G2997,G2991);
not gate_1008(G2998,G2994);
and gate_1009(G689,G681,G683);
and gate_1010(G700,G663,G694);
or gate_1011(G1539,G1536,G1537,G1538);
or gate_1012(G1584,G1582,G1583);
or gate_1013(G1588,G1586,G1587);
or gate_1014(G1592,G1590,G1591);
or gate_1015(G1596,G1594,G1595);
or gate_1016(G1600,G1598,G1599);
or gate_1017(G1604,G1602,G1603);
or gate_1018(G1608,G1606,G1607);
and gate_1019(G1661,G673,G1656);
or gate_1020(G1892,G1883,G1886);
nor gate_1021(G1893,G1883,G1886);
and gate_1022(G1933,G169,G1912,G1927);
and gate_1023(G1936,G179,G1912,G1930);
and gate_1024(G1939,G190,G1916,G1930);
and gate_1025(G1940,G200,G1916,G1927);
not gate_1026(G1941,G1916);
or gate_1027(G1993,G1984,G1987);
nor gate_1028(G1996,G1984,G1987);
or gate_1029(G2043,G2034,G2037);
nor gate_1030(G2046,G2034,G2037);
or gate_1031(G2100,G2091,G2094);
nor gate_1032(G2101,G2091,G2094);
and gate_1033(G2143,G169,G2120,G2137);
and gate_1034(G2146,G179,G2120,G2140);
and gate_1035(G2149,G190,G2124,G2140);
and gate_1036(G2150,G200,G2124,G2137);
not gate_1037(G2151,G2124);
or gate_1038(G2205,G2196,G2199);
nor gate_1039(G2208,G2196,G2199);
or gate_1040(G2257,G2248,G2251);
nor gate_1041(G2260,G2248,G2251);
not gate_1042(G3138,G3134);
and gate_1043(G2328,G2285,G1912);
not gate_1044(G3162,G3158);
not gate_1045(G3170,G3166);
not gate_1046(G3178,G3174);
not gate_1047(G3186,G3182);
not gate_1048(G3204,G3200);
and gate_1049(G2375,G2298,G2120);
not gate_1050(G3236,G3232);
not gate_1051(G3244,G3240);
not gate_1052(G3252,G3248);
not gate_1053(G3228,G3224);
buf gate_1054(G3066,G600);
buf gate_1055(G3074,G600);
not gate_1056(G3128,G3124);
not gate_1057(G3194,G3190);
nand gate_1058(G619,G2994,G2997);
nand gate_1059(G620,G2991,G2998);
nand gate_1060(G582,G3002,G3005);
nand gate_1061(G583,G2999,G3006);
or gate_1062(G692,G689,G690,G691);
or gate_1063(G703,G700,G701,G702);
and gate_1064(G1612,G1539,G1609);
and gate_1065(G1621,G1584,G1618);
and gate_1066(G1630,G1588,G1627);
and gate_1067(G1639,G1592,G1636);
and gate_1068(G1648,G1596,G1645);
and gate_1069(G1657,G1600,G1654);
and gate_1070(G1666,G1604,G1663);
and gate_1071(G1675,G1608,G1672);
and gate_1072(G1895,G1893,G1894);
or gate_1073(G1946,G1939,G1940,G1941);
and gate_1074(G1998,G1996,G1997);
and gate_1075(G2048,G2046,G2047);
and gate_1076(G2103,G2101,G2102);
or gate_1077(G2156,G2149,G2150,G2151);
and gate_1078(G2210,G2208,G2209);
and gate_1079(G2262,G2260,G2261);
not gate_1080(G2271,G1892);
not gate_1081(G2311,G2100);
nand gate_1082(G356,G619,G620);
nand gate_1083(G357,G582,G583);
nand gate_1084(G603,G3074,G3077);
not gate_1085(G3078,G3074);
nand gate_1086(G606,G3066,G3069);
not gate_1087(G3070,G3066);
and gate_1088(G1670,G703,G1665);
and gate_1089(G1679,G692,G1674);
or gate_1090(G1942,G1933,G1936);
nor gate_1091(G1945,G1933,G1936);
or gate_1092(G2152,G2143,G2146);
nor gate_1093(G2155,G2143,G2146);
and gate_1094(G2445,G1993,G2293);
and gate_1095(G2448,G2043,G2293);
and gate_1096(G2455,G2205,G2302);
and gate_1097(G2458,G2257,G2302);
buf gate_1098(G3142,G2328);
buf gate_1099(G3150,G2328);
buf gate_1100(G3208,G2375);
buf gate_1101(G3216,G2375);
nand gate_1102(G358,G356,G357);
nand gate_1103(G604,G3071,G3078);
nand gate_1104(G607,G3063,G3070);
and gate_1105(G1947,G1945,G1946);
and gate_1106(G2157,G2155,G2156);
buf gate_1107(G2317,G1895);
buf gate_1108(G2338,G1998);
buf gate_1109(G2351,G2048);
buf gate_1110(G2364,G2103);
buf gate_1111(G2380,G2210);
buf gate_1112(G2388,G2262);
nand gate_1113(G605,G603,G604);
nand gate_1114(G608,G606,G607);
nand gate_1115(G2272,G1895,G1942);
nand gate_1116(G2312,G2103,G2152);
not gate_1117(G3146,G3142);
not gate_1118(G3154,G3150);
not gate_1119(G3220,G3216);
not gate_1120(G3212,G3208);
and gate_1121(G2444,G1942,G2288);
buf gate_1122(G2451,G2448);
and gate_1123(G2454,G2152,G2293);
buf gate_1124(G2461,G2458);
not gate_1125(G2530,G2445);
buf gate_1126(G3323,G2458);
not gate_1127(G349,G605);
not gate_1128(G350,G608);
and gate_1129(G2265,G1895,G1947,G1998,G2048);
nand gate_1130(G2273,G1895,G1947,G1993);
nand gate_1131(G2274,G2043,G1947,G1998,G1895);
and gate_1132(G2309,G2103,G2157,G2210,G2262);
nand gate_1133(G2313,G2103,G2157,G2205);
nand gate_1134(G2314,G2257,G2157,G2210,G2103);
buf gate_1135(G2325,G1947);
buf gate_1136(G2372,G2157);
not gate_1137(G2523,G2444);
not gate_1138(G2533,G2454);
buf gate_1139(G3121,G2317);
buf gate_1140(G3131,G2317);
buf gate_1141(G3155,G2338);
buf gate_1142(G3163,G2338);
buf gate_1143(G3171,G2351);
buf gate_1144(G3179,G2351);
buf gate_1145(G3187,G2364);
buf gate_1146(G3197,G2364);
buf gate_1147(G3221,G2380);
buf gate_1148(G3229,G2380);
buf gate_1149(G3237,G2388);
buf gate_1150(G3245,G2388);
nand gate_1151(G351,G349,G350);
nand gate_1152(G2275,G2271,G2272,G2273,G2274);
nand gate_1153(G2315,G2311,G2312,G2313,G2314);
not gate_1154(G3329,G3323);
and gate_1155(G372,G2309,G2265);
nand gate_1156(G2324,G3131,G3138);
nand gate_1157(G2350,G3163,G3170);
nand gate_1158(G2363,G3179,G3186);
nand gate_1159(G2371,G3197,G3204);
nand gate_1160(G2387,G3229,G3236);
nand gate_1161(G2400,G3245,G3252);
buf gate_1162(G2268,G2265);
not gate_1163(G3137,G3131);
not gate_1164(G3161,G3155);
nand gate_1165(G2345,G3155,G3162);
not gate_1166(G3169,G3163);
not gate_1167(G3177,G3171);
nand gate_1168(G2358,G3171,G3178);
not gate_1169(G3185,G3179);
not gate_1170(G3203,G3197);
not gate_1171(G3235,G3229);
not gate_1172(G3243,G3237);
nand gate_1173(G2395,G3237,G3244);
not gate_1174(G3251,G3245);
not gate_1175(G3227,G3221);
nand gate_1176(G2432,G3221,G3228);
and gate_1177(G2490,G2309,G2485);
not gate_1178(G3127,G3121);
nand gate_1179(G3130,G3121,G3128);
buf gate_1180(G3139,G2325);
buf gate_1181(G3147,G2325);
not gate_1182(G3193,G3187);
nand gate_1183(G3196,G3187,G3194);
buf gate_1184(G3205,G2372);
buf gate_1185(G3213,G2372);
nand gate_1186(G2307,G2265,G2315);
not gate_1187(G2308,G2275);
nand gate_1188(G2323,G3134,G3137);
nand gate_1189(G2349,G3166,G3169);
nand gate_1190(G2362,G3182,G3185);
nand gate_1191(G2370,G3200,G3203);
nand gate_1192(G2386,G3232,G3235);
nand gate_1193(G2399,G3248,G3251);
nand gate_1194(G2344,G3158,G3161);
nand gate_1195(G2357,G3174,G3177);
nand gate_1196(G2394,G3240,G3243);
nand gate_1197(G2431,G3224,G3227);
and gate_1198(G2464,G2315,G2302);
or gate_1199(G2491,G2489,G2490);
nand gate_1200(G3129,G3124,G3127);
nand gate_1201(G3195,G3190,G3193);
and gate_1202(G368,G2307,G2308);
nand gate_1203(G1615,G2323,G2324);
nand gate_1204(G2337,G3147,G3154);
nand gate_1205(G1633,G2349,G2350);
nand gate_1206(G1642,G2362,G2363);
nand gate_1207(G1651,G2370,G2371);
nand gate_1208(G2379,G3213,G3220);
nand gate_1209(G1669,G2386,G2387);
nand gate_1210(G1678,G2399,G2400);
not gate_1211(G3145,G3139);
nand gate_1212(G2332,G3139,G3146);
not gate_1213(G3153,G3147);
nand gate_1214(G2346,G2344,G2345);
nand gate_1215(G2359,G2357,G2358);
not gate_1216(G3219,G3213);
nand gate_1217(G2396,G2394,G2395);
not gate_1218(G3211,G3205);
nand gate_1219(G2425,G3205,G3212);
nand gate_1220(G2433,G2431,G2432);
nand gate_1221(G3272,G3129,G3130);
nand gate_1222(G3308,G3195,G3196);
not gate_1223(G369,G368);
not gate_1224(G1613,G1615);
nand gate_1225(G2336,G3150,G3153);
not gate_1226(G1631,G1633);
not gate_1227(G1640,G1642);
not gate_1228(G1649,G1651);
nand gate_1229(G2378,G3216,G3219);
not gate_1230(G1667,G1669);
not gate_1231(G1676,G1678);
nand gate_1232(G2331,G3142,G3145);
nand gate_1233(G2424,G3208,G3211);
buf gate_1234(G2467,G2464);
buf gate_1235(G2495,G2491);
buf gate_1236(G3295,G2464);
and gate_1237(G3374,G330,G2491);
and gate_1238(G1614,G1613,G1610);
nand gate_1239(G1624,G2336,G2337);
and gate_1240(G1632,G1631,G1628);
and gate_1241(G1641,G1640,G1637);
and gate_1242(G1650,G1649,G1646);
nand gate_1243(G1660,G2378,G2379);
and gate_1244(G1668,G1667,G1664);
and gate_1245(G1677,G1676,G1673);
nand gate_1246(G2333,G2331,G2332);
buf gate_1247(G2406,G2346);
buf gate_1248(G2409,G2346);
buf gate_1249(G2415,G2359);
buf gate_1250(G2419,G2359);
nand gate_1251(G2426,G2424,G2425);
buf gate_1252(G2439,G2396);
and gate_1253(G2518,G2433,G2461);
not gate_1254(G3276,G3272);
not gate_1255(G3312,G3308);
and gate_1256(G2612,G330,G2396);
buf gate_1257(G3326,G2433);
nor gate_1258(G1617,G1612,G1614,G1616);
not gate_1259(G1622,G1624);
nor gate_1260(G1635,G1630,G1632,G1634);
nor gate_1261(G1644,G1639,G1641,G1643);
nor gate_1262(G1653,G1648,G1650,G1652);
not gate_1263(G1658,G1660);
nor gate_1264(G1671,G1666,G1668,G1670);
nor gate_1265(G1680,G1675,G1677,G1679);
and gate_1266(G2500,G2467,G2268);
and gate_1267(G2505,G2495,G2268);
or gate_1268(G2519,G2455,G2518);
not gate_1269(G3378,G3374);
not gate_1270(G2642,G2467);
buf gate_1271(G2645,G2467);
not gate_1272(G3301,G3295);
and gate_1273(G1623,G1622,G1619);
and gate_1274(G1659,G1658,G1655);
buf gate_1275(G2401,G2333);
or gate_1276(G2501,G2275,G2500);
and gate_1277(G2511,G2495,G2419,G2409);
and gate_1278(G2512,G2495,G2415);
and gate_1279(G2513,G2439,G2433,G2426);
and gate_1280(G2514,G2439,G2433);
and gate_1281(G2517,G2467,G2415);
nand gate_1282(G2531,G2409,G2451);
nand gate_1283(G2532,G2409,G2419,G2467);
nand gate_1284(G2534,G2426,G2455);
nand gate_1285(G2535,G2426,G2433,G2461);
nand gate_1286(G2607,G3326,G3329);
not gate_1287(G3330,G3326);
and gate_1288(G2643,G330,G2491,G2642);
and gate_1289(G2687,G1617,G2680);
and gate_1290(G2725,G1635,G2718);
and gate_1291(G2742,G1644,G2735);
and gate_1292(G2760,G1653,G2753);
and gate_1293(G2794,G1671,G2787);
and gate_1294(G2811,G1680,G2804);
buf gate_1295(G3280,G2333);
buf gate_1296(G3290,G2409);
buf gate_1297(G3298,G2415);
buf gate_1298(G3316,G2426);
buf gate_1299(G3406,G2612);
buf gate_1300(G3414,G2612);
and gate_1301(G3422,G2439,G2439);
nor gate_1302(G1626,G1621,G1623,G1625);
nor gate_1303(G1662,G1657,G1659,G1661);
and gate_1304(G2567,G330,G2512);
and gate_1305(G2589,G330,G2513);
nand gate_1306(G2608,G3323,G3330);
buf gate_1307(G2654,G2519);
buf gate_1308(G3253,G2505);
nand gate_1309(G3277,G2530,G2531,G2532);
or gate_1310(G3287,G2448,G2517);
nand gate_1311(G3305,G2533,G2534,G2535);
buf gate_1312(G3313,G2519);
and gate_1313(G3350,G330,G2511);
or gate_1314(G932,G2643,G2645);
and gate_1315(G2508,G2495,G2401,G2409,G2419);
nand gate_1316(G2524,G2401,G2445);
nand gate_1317(G2525,G2401,G2406,G2451);
nand gate_1318(G2526,G2401,G2406,G2419,G2467);
not gate_1319(G3294,G3290);
nand gate_1320(G2609,G2607,G2608);
not gate_1321(G3410,G3406);
not gate_1322(G3418,G3414);
nand gate_1323(G2624,G3422,G3425);
not gate_1324(G3426,G3422);
buf gate_1325(G2629,G2501);
nor gate_1326(G2647,G2643,G2645);
and gate_1327(G2706,G1626,G2699);
and gate_1328(G2777,G1662,G2770);
buf gate_1329(G3264,G2501);
not gate_1330(G3284,G3280);
not gate_1331(G3302,G3298);
nand gate_1332(G3303,G3298,G3301);
not gate_1333(G3320,G3316);
and gate_1334(G3398,G330,G2514);
not gate_1335(G2657,G2654);
and gate_1336(G398,G2519,G2654);
and gate_1337(G933,G932,G927);
nand gate_1338(G2527,G2523,G2524,G2525,G2526);
not gate_1339(G3259,G3253);
not gate_1340(G3354,G3350);
not gate_1341(G3293,G3287);
nand gate_1342(G2563,G3287,G3294);
not gate_1343(G3311,G3305);
nand gate_1344(G2585,G3305,G3312);
nand gate_1345(G2625,G3419,G3426);
not gate_1346(G3283,G3277);
nand gate_1347(G3286,G3277,G3284);
nand gate_1348(G3304,G3295,G3302);
not gate_1349(G3319,G3313);
nand gate_1350(G3322,G3313,G3320);
buf gate_1351(G3358,G2567);
buf gate_1352(G3366,G2567);
buf gate_1353(G3382,G2589);
buf gate_1354(G3390,G2589);
and gate_1355(G397,G330,G2514,G2657);
and gate_1356(G2544,G330,G2508);
nand gate_1357(G2562,G3290,G3293);
nand gate_1358(G2584,G3308,G3311);
not gate_1359(G3402,G3398);
nand gate_1360(G2626,G2624,G2625);
not gate_1361(G2632,G2629);
and gate_1362(G2634,G2501,G2629);
buf gate_1363(G2650,G2647);
not gate_1364(G3268,G3264);
buf gate_1365(G3256,G2508);
nand gate_1366(G3285,G3280,G3283);
nand gate_1367(G3321,G3316,G3319);
nand gate_1368(G3371,G3303,G3304);
buf gate_1369(G3403,G2609);
buf gate_1370(G3411,G2609);
or gate_1371(G362,G929,G933,G938);
nor gate_1372(G1030,G929,G933,G938);
or gate_1373(G399,G397,G398);
nand gate_1374(G2564,G2562,G2563);
not gate_1375(G3362,G3358);
not gate_1376(G3370,G3366);
nand gate_1377(G2586,G2584,G2585);
not gate_1378(G3386,G3382);
not gate_1379(G3394,G3390);
and gate_1380(G2633,G330,G2505,G2632);
buf gate_1381(G3261,G2527);
buf gate_1382(G3269,G2527);
nand gate_1383(G3347,G3285,G3286);
nand gate_1384(G3395,G3321,G3322);
not gate_1385(G363,G1030);
nand gate_1386(G2536,G3256,G3259);
not gate_1387(G3260,G3256);
not gate_1388(G3377,G3371);
nand gate_1389(G2580,G3371,G3378);
not gate_1390(G3409,G3403);
nand gate_1391(G2616,G3403,G3410);
not gate_1392(G3417,G3411);
nand gate_1393(G2622,G3411,G3418);
nor gate_1394(G2635,G2633,G2634);
and gate_1395(G2805,G2626,G2802);
and gate_1396(G2808,G2626,G2803);
buf gate_1397(G3334,G2544);
buf gate_1398(G3342,G2544);
buf gate_1399(G3454,G2650);
and gate_1400(G364,G362,G363);
nand gate_1401(G2537,G3253,G3260);
not gate_1402(G3275,G3269);
nand gate_1403(G2540,G3269,G3276);
not gate_1404(G3353,G3347);
nand gate_1405(G2557,G3347,G3354);
nand gate_1406(G2579,G3374,G3377);
not gate_1407(G3401,G3395);
nand gate_1408(G2602,G3395,G3402);
nand gate_1409(G2615,G3406,G3409);
nand gate_1410(G2621,G3414,G3417);
not gate_1411(G3267,G3261);
nand gate_1412(G3112,G3261,G3268);
buf gate_1413(G3355,G2564);
buf gate_1414(G3363,G2564);
buf gate_1415(G3379,G2586);
buf gate_1416(G3387,G2586);
nand gate_1417(G2538,G2536,G2537);
nand gate_1418(G2539,G3272,G3275);
not gate_1419(G3338,G3334);
not gate_1420(G3346,G3342);
nand gate_1421(G2556,G3350,G3353);
nand gate_1422(G2581,G2579,G2580);
nand gate_1423(G2601,G3398,G3401);
nand gate_1424(G2617,G2615,G2616);
nand gate_1425(G2623,G2621,G2622);
buf gate_1426(G2638,G2635);
not gate_1427(G3458,G3454);
or gate_1428(G2814,G2805,G2808,G2811);
nor gate_1429(G2816,G2805,G2808,G2811);
nand gate_1430(G3111,G3264,G3267);
nand gate_1431(G2541,G2539,G2540);
nand gate_1432(G2558,G2556,G2557);
not gate_1433(G3361,G3355);
nand gate_1434(G2571,G3355,G3362);
not gate_1435(G3369,G3363);
nand gate_1436(G2577,G3363,G3370);
not gate_1437(G3385,G3379);
nand gate_1438(G2593,G3379,G3386);
not gate_1439(G3393,G3387);
nand gate_1440(G2598,G3387,G3394);
nand gate_1441(G2603,G2601,G2602);
nand gate_1442(G3113,G3111,G3112);
and gate_1443(G3116,G330,G2538);
not gate_1444(G3451,G2623);
not gate_1445(G395,G2816);
nand gate_1446(G2570,G3358,G3361);
nand gate_1447(G2576,G3366,G3369);
nand gate_1448(G2592,G3382,G3385);
nand gate_1449(G2597,G3390,G3393);
and gate_1450(G2736,G2581,G2733);
and gate_1451(G2739,G2581,G2734);
and gate_1452(G2788,G2617,G2785);
buf gate_1453(G3438,G2638);
and gate_1454(G3446,G2617,G2647);
buf gate_1455(G3459,G2814);
and gate_1456(G396,G2814,G395);
not gate_1457(G3119,G3113);
not gate_1458(G3120,G3116);
nand gate_1459(G2572,G2570,G2571);
nand gate_1460(G2578,G2576,G2577);
nand gate_1461(G2594,G2592,G2593);
nand gate_1462(G2599,G2597,G2598);
nand gate_1463(G2677,G3451,G3458);
not gate_1464(G3457,G3451);
and gate_1465(G2700,G2558,G2697);
and gate_1466(G2771,G2603,G2768);
buf gate_1467(G3331,G2541);
buf gate_1468(G3339,G2541);
buf gate_1469(G3427,G2558);
buf gate_1470(G3443,G2603);
nand gate_1471(G954,G3116,G3119);
nand gate_1472(G955,G3113,G3120);
not gate_1473(G2600,G2599);
not gate_1474(G3442,G3438);
not gate_1475(G3450,G3446);
nand gate_1476(G2676,G3454,G3457);
or gate_1477(G2745,G2736,G2739,G2742);
nor gate_1478(G2748,G2736,G2739,G2742);
not gate_1479(G3465,G3459);
not gate_1480(G3435,G2578);
nand gate_1481(G950,G954,G955);
not gate_1482(G3337,G3331);
nand gate_1483(G2548,G3331,G3338);
not gate_1484(G3345,G3339);
nand gate_1485(G2553,G3339,G3346);
nor gate_1486(G2661,G2600,G2650);
and gate_1487(G2662,G2617,G2603,G2594,G2650);
not gate_1488(G3433,G3427);
not gate_1489(G3449,G3443);
nand gate_1490(G2672,G3443,G3450);
nand gate_1491(G2674,G2676,G2677);
and gate_1492(G2719,G2572,G2716);
and gate_1493(G2754,G2594,G2751);
and gate_1494(G3430,G2572,G2635);
not gate_1495(G383,G2748);
and gate_1496(G951,G950,G943);
nand gate_1497(G2547,G3334,G3337);
nand gate_1498(G2552,G3342,G3345);
or gate_1499(G2663,G2661,G2662);
nand gate_1500(G2670,G3435,G3442);
not gate_1501(G3441,G3435);
nand gate_1502(G2671,G3446,G3449);
not gate_1503(G2675,G2674);
buf gate_1504(G3491,G2745);
buf gate_1505(G3499,G2745);
and gate_1506(G384,G2745,G383);
nand gate_1507(G2549,G2547,G2548);
nand gate_1508(G2554,G2552,G2553);
nand gate_1509(G2664,G3430,G3433);
not gate_1510(G3434,G3430);
nand gate_1511(G2669,G3438,G3441);
nand gate_1512(G2673,G2671,G2672);
and gate_1513(G2757,G2663,G2752);
and gate_1514(G2791,G2675,G2786);
or gate_1515(G365,G944,G947,G951);
nor gate_1516(G1031,G944,G947,G951);
not gate_1517(G2555,G2554);
nand gate_1518(G2665,G3427,G3434);
nand gate_1519(G2667,G2669,G2670);
and gate_1520(G2774,G2673,G2769);
not gate_1521(G3497,G3491);
not gate_1522(G3505,G3499);
not gate_1523(G366,G1031);
nor gate_1524(G2658,G2555,G2638);
and gate_1525(G2659,G2572,G2558,G2549,G2638);
nand gate_1526(G2666,G2664,G2665);
not gate_1527(G2668,G2667);
and gate_1528(G2681,G2549,G2678);
or gate_1529(G2763,G2754,G2757,G2760);
nor gate_1530(G2765,G2754,G2757,G2760);
or gate_1531(G2797,G2788,G2791,G2794);
nor gate_1532(G2799,G2788,G2791,G2794);
and gate_1533(G367,G365,G366);
or gate_1534(G2660,G2658,G2659);
and gate_1535(G2703,G2666,G2698);
and gate_1536(G2722,G2668,G2717);
or gate_1537(G2780,G2771,G2774,G2777);
nor gate_1538(G2782,G2771,G2774,G2777);
not gate_1539(G386,G2765);
not gate_1540(G392,G2799);
and gate_1541(G2684,G2660,G2679);
buf gate_1542(G3462,G2797);
buf gate_1543(G3470,G2763);
and gate_1544(G387,G2763,G386);
not gate_1545(G389,G2782);
and gate_1546(G393,G2797,G392);
or gate_1547(G2709,G2700,G2703,G2706);
nor gate_1548(G2713,G2700,G2703,G2706);
or gate_1549(G2728,G2719,G2722,G2725);
nor gate_1550(G2730,G2719,G2722,G2725);
and gate_1551(G2922,G2816,G2799,G2782,G2765);
buf gate_1552(G3467,G2780);
and gate_1553(G390,G2780,G389);
or gate_1554(G2690,G2681,G2684,G2687);
nor gate_1555(G2694,G2681,G2684,G2687);
nand gate_1556(G2821,G3462,G3465);
not gate_1557(G3466,G3462);
not gate_1558(G3474,G3470);
and gate_1559(G378,G2709,G2709);
not gate_1560(G380,G2730);
nand gate_1561(G2822,G3459,G3466);
not gate_1562(G3473,G3467);
nand gate_1563(G2827,G3467,G3474);
buf gate_1564(G2839,G2728);
and gate_1565(G2883,G2709,G2871);
buf gate_1566(G3507,G2709);
and gate_1567(G375,G2690,G2690);
and gate_1568(G381,G2728,G380);
nand gate_1569(G2823,G2821,G2822);
nand gate_1570(G2826,G3470,G3473);
and gate_1571(G2880,G2871,G2690);
and gate_1572(G2925,G2748,G2730,G2713,G2694);
and gate_1573(G2928,G2713,G2694,G2874);
buf gate_1574(G3510,G2690);
nand gate_1575(G2828,G2826,G2827);
buf gate_1576(G3494,G2839);
buf gate_1577(G3502,G2839);
not gate_1578(G3513,G3507);
buf gate_1579(G3544,G2883);
buf gate_1580(G3552,G2883);
and gate_1581(G406,G2922,G2925);
and gate_1582(G2929,G2922,G2925);
buf gate_1583(G3475,G2823);
buf gate_1584(G3483,G2823);
not gate_1585(G3514,G3510);
nand gate_1586(G3515,G3510,G3513);
buf gate_1587(G3541,G2880);
buf gate_1588(G3549,G2880);
not gate_1589(G407,G406);
nor gate_1590(G2930,G2928,G2929);
nand gate_1591(G2842,G3494,G3497);
not gate_1592(G3498,G3494);
nand gate_1593(G2852,G3502,G3505);
not gate_1594(G3506,G3502);
not gate_1595(G3548,G3544);
not gate_1596(G3556,G3552);
buf gate_1597(G3478,G2828);
buf gate_1598(G3486,G2828);
nand gate_1599(G3516,G3507,G3514);
and gate_1600(G408,G213,G2930);
not gate_1601(G3481,G3475);
not gate_1602(G3489,G3483);
nand gate_1603(G2843,G3491,G3498);
nand gate_1604(G2853,G3499,G3506);
not gate_1605(G3547,G3541);
nand gate_1606(G2887,G3541,G3548);
nand gate_1607(G2896,G3549,G3556);
not gate_1608(G3555,G3549);
nand gate_1609(G3520,G3515,G3516);
not gate_1610(G409,G408);
nand gate_1611(G2831,G3478,G3481);
not gate_1612(G3482,G3478);
nand gate_1613(G2836,G3486,G3489);
not gate_1614(G3490,G3486);
nand gate_1615(G2844,G2842,G2843);
nand gate_1616(G2848,G2852,G2853);
nand gate_1617(G2886,G3544,G3547);
nand gate_1618(G2895,G3552,G3555);
nand gate_1619(G2832,G3475,G3482);
nand gate_1620(G2837,G3483,G3490);
not gate_1621(G2849,G2848);
not gate_1622(G3524,G3520);
nand gate_1623(G2888,G2886,G2887);
nand gate_1624(G2891,G2895,G2896);
nand gate_1625(G2833,G2831,G2832);
nand gate_1626(G2838,G2836,G2837);
not gate_1627(G2892,G2891);
buf gate_1628(G3517,G2844);
and gate_1629(G2906,G2844,G2888,G2900);
and gate_1630(G2908,G2849,G2888,G2903);
not gate_1631(G2913,G2838);
not gate_1632(G3523,G3517);
nand gate_1633(G2855,G3517,G3524);
and gate_1634(G2907,G2844,G2892,G2903);
and gate_1635(G2909,G2849,G2892,G2900);
buf gate_1636(G3525,G2833);
buf gate_1637(G3533,G2833);
nand gate_1638(G2854,G3520,G3523);
or gate_1639(G2910,G2906,G2907,G2908,G2909);
buf gate_1640(G3560,G2913);
buf gate_1641(G3568,G2913);
nand gate_1642(G2856,G2854,G2855);
not gate_1643(G3539,G3533);
not gate_1644(G3531,G3525);
not gate_1645(G3572,G3568);
not gate_1646(G3564,G3560);
buf gate_1647(G3557,G2910);
buf gate_1648(G3565,G2910);
buf gate_1649(G3528,G2856);
buf gate_1650(G3536,G2856);
nand gate_1651(G2921,G3557,G3564);
nand gate_1652(G2917,G3565,G3572);
not gate_1653(G3571,G3565);
not gate_1654(G3563,G3557);
nand gate_1655(G2863,G3528,G3531);
nand gate_1656(G2859,G3536,G3539);
nand gate_1657(G2920,G3560,G3563);
nand gate_1658(G2916,G3568,G3571);
not gate_1659(G3540,G3536);
not gate_1660(G3532,G3528);
nand gate_1661(G2864,G3525,G3532);
nand gate_1662(G2860,G3533,G3540);
nand gate_1663(G403,G2920,G2921);
nand gate_1664(G404,G2916,G2917);
nand gate_1665(G400,G2863,G2864);
nand gate_1666(G401,G2859,G2860);
and gate_1667(G405,G403,G404);
nand gate_1668(G402,G400,G401);
endmodule
