module test(a, c);
    input wire a;
    output wire [3:0] c;
    assign c = 4'b0001;

endmodule
