// Verilog File 
module c2670 (G1,G2,G3,G4,G5,G6,G7,G8,G11,
G14,G15,G16,G19,G20,G21,G22,G23,G24,G25,
G26,G27,G28,G29,G32,G33,G34,G35,G36,G37,
G40,G43,G44,G47,G48,G49,G50,G51,G52,G53,
G54,G55,G56,G57,G60,G61,G62,G63,G64,G65,
G66,G67,G68,G69,G72,G73,G74,G75,G76,G77,
G78,G79,G80,G81,G82,G85,G86,G87,G88,G89,
G90,G91,G92,G93,G94,G95,G96,G99,G100,G101,
G102,G103,G104,G105,G106,G107,G108,G111,G112,G113,
G114,G115,G116,G117,G118,G119,G120,G123,G124,G125,
G126,G127,G128,G129,G130,G131,G132,G135,G136,G137,
G138,G139,G140,G141,G142,G452,G483,G543,G559,G567,
G651,G661,G860,G868,G1083,G1341,G1348,G1384,G1956,G1961,
G1966,G1971,G1976,G1981,G1986,G1991,G1996,G2066,G2067,G2072,
G2078,G2084,G2090,G2096,G2100,G2104,G2105,G2106,G2427,G2430,
G2435,G2438,G2443,G2446,G2451,G2454,G2474,G2678,G350,G335,
G409,G369,G367,G411,G337,G384,G218,G219,G220,G221,
G235,G236,G237,G238,G158,G259,G391,G173,G223,G234,
G217,G325,G261,G319,G160,G162,G164,G166,G168,G171,
G153,G176,G188,G299,G301,G286,G303,G288,G305,G290,
G284,G321,G297,G280,G148,G282,G323,G156,G401,G227,
G229,G311,G150,G145,G395,G295,G331,G397,G329,G231,
G308,G225);

input G1,G2,G3,G4,G5,G6,G7,G8,G11,
G14,G15,G16,G19,G20,G21,G22,G23,G24,G25,
G26,G27,G28,G29,G32,G33,G34,G35,G36,G37,
G40,G43,G44,G47,G48,G49,G50,G51,G52,G53,
G54,G55,G56,G57,G60,G61,G62,G63,G64,G65,
G66,G67,G68,G69,G72,G73,G74,G75,G76,G77,
G78,G79,G80,G81,G82,G85,G86,G87,G88,G89,
G90,G91,G92,G93,G94,G95,G96,G99,G100,G101,
G102,G103,G104,G105,G106,G107,G108,G111,G112,G113,
G114,G115,G116,G117,G118,G119,G120,G123,G124,G125,
G126,G127,G128,G129,G130,G131,G132,G135,G136,G137,
G138,G139,G140,G141,G142,G452,G483,G543,G559,G567,
G651,G661,G860,G868,G1083,G1341,G1348,G1384,G1956,G1961,
G1966,G1971,G1976,G1981,G1986,G1991,G1996,G2066,G2067,G2072,
G2078,G2084,G2090,G2096,G2100,G2104,G2105,G2106,G2427,G2430,
G2435,G2438,G2443,G2446,G2451,G2454,G2474,G2678;

output G350,G335,G409,G369,G367,G411,G337,G384,G218,
G219,G220,G221,G235,G236,G237,G238,G158,G259,G391,
G173,G223,G234,G217,G325,G261,G319,G160,G162,G164,
G166,G168,G171,G153,G176,G188,G299,G301,G286,G303,
G288,G305,G290,G284,G321,G297,G280,G148,G282,G323,
G156,G401,G227,G229,G311,G150,G145,G395,G295,G331,
G397,G329,G231,G308,G225;

wire G546,G560,G1385,G157,G547,G258,G480,G486,G654,
G655,G658,G772,G795,G865,G875,G882,G1251,G1254,G1261,
G1284,G1344,G1351,G1394,G1418,G2433,G2434,G2441,G2442,G2449,
G2450,G2478,G1631,G1655,G1710,G1721,G2682,G1955,G1959,G1964,
G1969,G1974,G1979,G1984,G1989,G1994,G1999,G2001,G2012,G2070,
G2076,G2082,G2088,G2094,G2099,G2103,G2457,G2458,G2461,G2464,
G2471,G2479,G2482,G2487,G2490,G2495,G2498,G2505,G2508,G2675,
G2683,G2686,G2691,G2694,G2699,G2702,G487,G1475,G1476,G1484,
G1485,G1493,G1494,G2459,G2460,G216,G1253,G1256,G558,G748,
G784,G807,G821,G825,G829,G833,G837,G881,G994,G1273,
G1296,G1310,G1314,G1318,G1322,G1326,G1406,G1430,G1444,G1448,
G1452,G1456,G1460,G1477,G1486,G1495,G2477,G1499,G2485,G2486,
G2493,G2494,G1643,G1667,G1681,G1685,G1689,G1693,G1697,G1716,
G1728,G2681,G1776,G2689,G2690,G2697,G2698,G1831,G1893,G2007,
G2018,G2467,G2468,G2501,G2502,G2511,G2512,G2518,G2551,G2559,
G2567,G2575,G2583,G2591,G2599,G2607,G2615,G2623,G2705,G2706,
G2735,G2743,G2751,G2759,G2767,G2775,G550,G552,G894,G1498,
G1507,G1508,G1516,G1517,G1775,G1784,G1785,G1793,G1794,G2469,
G2470,G2503,G2504,G2513,G2514,G2707,G2708,G551,G553,G818,
G819,G820,G822,G823,G824,G826,G827,G828,G830,G831,
G832,G834,G835,G836,G1307,G1308,G1309,G1311,G1312,G1313,
G1315,G1316,G1317,G1319,G1320,G1321,G1323,G1324,G1325,G1441,
G1442,G1443,G1445,G1446,G1447,G1449,G1450,G1451,G1453,G1454,
G1455,G1457,G1458,G1459,G1481,G1490,G1500,G1509,G1518,G1521,
G1525,G2557,G2565,G2573,G2581,G2589,G2597,G2605,G2613,G2621,
G2629,G1678,G1679,G1680,G1682,G1683,G1684,G1686,G1687,G1688,
G1690,G1691,G1692,G1694,G1695,G1696,G1734,G1736,G1738,G1740,
G1742,G1744,G1746,G1748,G1750,G1777,G1786,G1795,G2023,G2025,
G2027,G2029,G2031,G2033,G2035,G2037,G2741,G2749,G2757,G2765,
G2773,G2781,G2515,G2522,G2525,G2528,G2730,G554,G838,G841,
G846,G854,G857,G1327,G1329,G1331,G1333,G1335,G1461,G1464,
G1467,G1470,G1473,G1698,G1701,G1704,G1707,G2634,G1504,G1513,
G1524,G1528,G1529,G1533,G1538,G1541,G1781,G1790,G1806,G1810,
G2734,G2521,G2524,G2531,G2532,G144,G147,G152,G175,G187,
G516,G852,G885,G887,G893,G1028,G1031,G1035,G1041,G1049,
G1057,G1060,G1066,G1072,G1078,G1213,G1218,G1250,G1387,G1389,
G1537,G1540,G1735,G1737,G1739,G1741,G1743,G1745,G1747,G1749,
G1751,G2638,G2024,G2026,G2028,G2030,G2032,G2034,G2036,G2038,
G2154,G2523,G2533,G2534,G2631,G2639,G2642,G2647,G2650,G2655,
G2658,G2665,G2668,G1532,G1536,G1539,G1542,G1544,G1547,G2065,
G1809,G1813,G1821,G1824,G2538,G2546,G2554,G2562,G2570,G2578,
G2586,G2594,G2602,G2610,G2618,G2626,G2738,G2746,G2754,G2762,
G2770,G2778,G456,G466,G562,G883,G889,G891,G1043,G1051,
G1062,G1068,G1074,G1080,G1225,G1227,G1232,G1234,G1543,G1546,
G2637,G1753,G2645,G2646,G2653,G2654,G1820,G1823,G2107,G2110,
G2118,G2123,G2151,G2158,G2161,G2164,G2172,G2235,G2262,G2350,
G2535,G2661,G2662,G2671,G2672,G468,G897,G898,G1228,G1235,
G1545,G1548,G2542,G2550,G1561,G2558,G1565,G2566,G1569,G2574,
G1573,G2582,G1577,G2590,G1581,G2598,G1585,G2606,G1589,G2614,
G1593,G2622,G1597,G2630,G1752,G1761,G1762,G1770,G1771,G1822,
G1825,G2039,G2742,G2043,G2750,G2047,G2758,G2051,G2766,G2055,
G2774,G2059,G2782,G2663,G2664,G2673,G2674,G146,G462,G2113,
G2114,G2122,G2129,G592,G2167,G2168,G2176,G2241,G2266,G743,
G749,G886,G995,G1006,G1550,G2354,G2541,G1562,G1566,G1570,
G1574,G1578,G1582,G1586,G1590,G1594,G1598,G1754,G1763,G1772,
G2040,G2044,G2048,G2052,G2056,G2060,G2115,G2126,G2131,G2134,
G2141,G2144,G2157,G2160,G2169,G2177,G2180,G2187,G2190,G2207,
G2254,G2334,G2342,G2422,G2543,G2709,G2712,G2727,G569,G570,
G599,G600,G896,G1549,G1243,G1245,G1257,G1258,G1563,G1567,
G1571,G1575,G1579,G1583,G1587,G1591,G1595,G1599,G2041,G2045,
G2049,G2053,G2057,G2061,G2159,G475,G490,G496,G502,G508,
G765,G769,G571,G2121,G579,G587,G2130,G596,G601,G2175,
G609,G2258,G1014,G1018,G717,G723,G729,G735,G753,G2338,
G999,G1091,G2346,G2426,G1337,G2549,G1552,G1600,G1596,G1592,
G1588,G1584,G1580,G1576,G1572,G1568,G1564,G2062,G2058,G2054,
G2050,G2046,G2042,G1758,G1767,G1798,G1802,G2733,G1829,G2137,
G2138,G2147,G2148,G2183,G2184,G2193,G2194,G2210,G2213,G2715,
G2716,G1094,G1096,G578,G588,G608,G742,G1005,G1092,G1551,
G1554,G1555,G1557,G1558,G1828,G1845,G1907,G2139,G2140,G2149,
G2150,G2185,G2186,G2195,G2196,G2717,G2718,G154,G155,G763,
G767,G531,G537,G575,G580,G589,G605,G610,G1012,G1016,
G705,G711,G1093,G1355,G1553,G1556,G1559,G1601,G1801,G1805,
G1815,G1818,G1830,G1836,G1850,G1898,G1912,G2197,G2200,G2214,
G2215,G2217,G2220,G2722,G492,G498,G504,G510,G519,G525,
G533,G539,G693,G699,G707,G713,G719,G725,G731,G737,
G1560,G1814,G1817,G2216,G493,G499,G505,G511,G521,G527,
G534,G540,G584,G613,G617,G621,G625,G676,G695,G701,
G708,G714,G720,G726,G732,G738,G1087,G1108,G1361,G1369,
G1373,G1377,G1607,G1615,G1619,G1623,G1816,G1819,G2726,G1842,
G1858,G1863,G1866,G1868,G1870,G1872,G1874,G1876,G1904,G1920,
G1925,G1928,G1930,G1932,G1934,G1936,G1938,G2203,G2204,G2223,
G2224,G2238,G522,G528,G696,G702,G1881,G1883,G1885,G1887,
G1889,G1891,G1943,G1945,G1947,G1949,G1951,G1953,G2205,G2206,
G2225,G2226,G2719,G616,G620,G624,G628,G630,G633,G636,
G639,G645,G2242,G675,G1107,G1368,G1371,G1375,G1614,G1617,
G1621,G1856,G1861,G1918,G1923,G2230,G2246,G2270,G2278,G2286,
G2294,G2302,G2310,G2358,G2366,G2374,G2382,G2390,G2398,G629,
G632,G635,G638,G646,G677,G1827,G907,G915,G922,G924,
G937,G946,G1109,G1125,G1133,G1140,G1142,G1155,G1164,G1378,
G1380,G1382,G1624,G1626,G1628,G2725,G1859,G1864,G1921,G1926,
G2267,G2275,G2283,G2291,G2299,G2307,G2318,G2326,G2355,G2363,
G2371,G2379,G2387,G2395,G2406,G2414,G647,G631,G634,G637,
G640,G2234,G2250,G679,G1826,G2274,G2282,G2290,G2298,G2306,
G2314,G1110,G2362,G2370,G2378,G2386,G2394,G2402,G1877,G1879,
G1939,G1941,G143,G671,G674,G686,G2273,G900,G2281,G909,
G2289,G917,G2297,G926,G2305,G929,G2313,G939,G2322,G2330,
G967,G1104,G1106,G2361,G1118,G2369,G1127,G2377,G1135,G2385,
G1144,G2393,G1147,G2401,G1157,G2410,G2418,G1184,G2227,G2243,
G2251,G2259,G2331,G2339,G2347,G2419,G687,G899,G908,G916,
G925,G928,G938,G954,G961,G1117,G1126,G1134,G1143,G1146,
G1156,G1172,G1179,G2315,G2323,G2403,G2411,G2233,G642,G2249,
G649,G2257,G665,G684,G2265,G688,G901,G910,G918,G927,
G930,G940,G2337,G963,G2345,G1099,G1115,G2353,G1119,G1128,
G1136,G1145,G1148,G1158,G2425,G1181,G641,G648,G664,G683,
G2321,G948,G2329,G956,G962,G1098,G1114,G2409,G1166,G2417,
G1174,G1180,G643,G650,G666,G681,G690,G947,G955,G964,
G968,G970,G971,G972,G978,G979,G1100,G1112,G1165,G1173,
G1182,G1185,G1187,G1188,G1189,G1195,G1196,G644,G884,G949,
G957,G969,G973,G1167,G1175,G1186,G1190,G680,G682,G895,
G1025,G1111,G1113,G685,G976,G977,G980,G981,G1116,G1193,
G1194,G1197,G1198,G982,G983,G988,G1027,G1199,G1200,G1205,
G984,G1085,G1201,G987,G990,G1204,G1207,G989,G1206,G991,
G1208,G1221,G1238,G1239,G1240,G1247,G471,G473,G1088,G1089;
buf gate_0(G350,G452);
buf gate_1(G335,G452);
buf gate_2(G409,G452);
and gate_3(G546,G1,G3);
not gate_4(G560,G559);
buf gate_5(G369,G1083);
buf gate_6(G367,G1083);
not gate_7(G1385,G1384);
buf gate_8(G411,G2066);
buf gate_9(G337,G2066);
buf gate_10(G384,G2066);
and gate_11(G157,G2090,G2084,G2078,G2072);
not gate_12(G547,G546);
not gate_13(G218,G44);
not gate_14(G219,G132);
not gate_15(G220,G82);
not gate_16(G221,G96);
not gate_17(G235,G69);
not gate_18(G236,G120);
not gate_19(G237,G57);
not gate_20(G238,G108);
and gate_21(G258,G2,G15,G661);
buf gate_22(G480,G661);
and gate_23(G486,G37,G37);
buf gate_24(G654,G452);
buf gate_25(G655,G8);
buf gate_26(G658,G8);
buf gate_27(G772,G543);
buf gate_28(G795,G651);
not gate_29(G865,G860);
not gate_30(G875,G868);
and gate_31(G882,G11,G868);
and gate_32(G1251,G132,G82,G96,G44);
and gate_33(G1254,G120,G57,G108,G69);
buf gate_34(G1261,G543);
buf gate_35(G1284,G651);
not gate_36(G1344,G1341);
not gate_37(G1351,G1348);
buf gate_38(G1394,G2104);
buf gate_39(G1418,G2105);
not gate_40(G2433,G2427);
not gate_41(G2434,G2430);
not gate_42(G2441,G2435);
not gate_43(G2442,G2438);
not gate_44(G2449,G2443);
not gate_45(G2450,G2446);
not gate_46(G2478,G2474);
buf gate_47(G1631,G2104);
buf gate_48(G1655,G2105);
buf gate_49(G1710,G16);
buf gate_50(G1721,G16);
not gate_51(G2682,G2678);
and gate_52(G1955,G7,G661);
not gate_53(G1959,G1956);
not gate_54(G1964,G1961);
not gate_55(G1969,G1966);
not gate_56(G1974,G1971);
not gate_57(G1979,G1976);
not gate_58(G1984,G1981);
not gate_59(G1989,G1986);
not gate_60(G1994,G1991);
not gate_61(G1999,G1996);
buf gate_62(G2001,G29);
buf gate_63(G2012,G29);
not gate_64(G2070,G2067);
not gate_65(G2076,G2072);
not gate_66(G2082,G2078);
not gate_67(G2088,G2084);
not gate_68(G2094,G2090);
not gate_69(G2099,G2096);
not gate_70(G2103,G2100);
not gate_71(G2457,G2451);
not gate_72(G2458,G2454);
buf gate_73(G2461,G1348);
buf gate_74(G2464,G1341);
buf gate_75(G2471,G1956);
buf gate_76(G2479,G1966);
buf gate_77(G2482,G1961);
buf gate_78(G2487,G1976);
buf gate_79(G2490,G1971);
buf gate_80(G2495,G1986);
buf gate_81(G2498,G1981);
buf gate_82(G2505,G1996);
buf gate_83(G2508,G1991);
buf gate_84(G2675,G2067);
buf gate_85(G2683,G2078);
buf gate_86(G2686,G2072);
buf gate_87(G2691,G2090);
buf gate_88(G2694,G2084);
buf gate_89(G2699,G2100);
buf gate_90(G2702,G2096);
not gate_91(G158,G157);
not gate_92(G259,G258);
not gate_93(G487,G486);
buf gate_94(G391,G654);
nand gate_95(G1475,G2430,G2433);
nand gate_96(G1476,G2427,G2434);
nand gate_97(G1484,G2438,G2441);
nand gate_98(G1485,G2435,G2442);
nand gate_99(G1493,G2446,G2449);
nand gate_100(G1494,G2443,G2450);
nand gate_101(G2459,G2454,G2457);
nand gate_102(G2460,G2451,G2458);
and gate_103(G173,G94,G654);
and gate_104(G216,G2106,G1955);
not gate_105(G223,G1955);
nand gate_106(G234,G567,G1955);
not gate_107(G1253,G1251);
not gate_108(G1256,G1254);
and gate_109(G558,G1254,G1251);
buf gate_110(G748,G655);
not gate_111(G784,G772);
not gate_112(G807,G795);
and gate_113(G821,G80,G772,G795);
and gate_114(G825,G68,G772,G795);
and gate_115(G829,G79,G772,G795);
and gate_116(G833,G78,G772,G795);
and gate_117(G837,G77,G772,G795);
and gate_118(G881,G11,G875);
buf gate_119(G994,G655);
not gate_120(G1273,G1261);
not gate_121(G1296,G1284);
and gate_122(G1310,G76,G1261,G1284);
and gate_123(G1314,G75,G1261,G1284);
and gate_124(G1318,G74,G1261,G1284);
and gate_125(G1322,G73,G1261,G1284);
and gate_126(G1326,G72,G1261,G1284);
not gate_127(G1406,G1394);
not gate_128(G1430,G1418);
and gate_129(G1444,G114,G1394,G1418);
and gate_130(G1448,G113,G1394,G1418);
and gate_131(G1452,G112,G1394,G1418);
and gate_132(G1456,G111,G1394,G1418);
and gate_133(G1460,G1394,G1418);
nand gate_134(G1477,G1475,G1476);
nand gate_135(G1486,G1484,G1485);
nand gate_136(G1495,G1493,G1494);
not gate_137(G2477,G2471);
nand gate_138(G1499,G2471,G2478);
not gate_139(G2485,G2479);
not gate_140(G2486,G2482);
not gate_141(G2493,G2487);
not gate_142(G2494,G2490);
not gate_143(G1643,G1631);
not gate_144(G1667,G1655);
and gate_145(G1681,G118,G1631,G1655);
and gate_146(G1685,G107,G1631,G1655);
and gate_147(G1689,G117,G1631,G1655);
and gate_148(G1693,G116,G1631,G1655);
and gate_149(G1697,G115,G1631,G1655);
not gate_150(G1716,G1710);
not gate_151(G1728,G1721);
not gate_152(G2681,G2675);
nand gate_153(G1776,G2675,G2682);
not gate_154(G2689,G2683);
not gate_155(G2690,G2686);
not gate_156(G2697,G2691);
not gate_157(G2698,G2694);
buf gate_158(G1831,G658);
buf gate_159(G1893,G658);
not gate_160(G2007,G2001);
not gate_161(G2018,G2012);
not gate_162(G2467,G2461);
not gate_163(G2468,G2464);
not gate_164(G2501,G2495);
not gate_165(G2502,G2498);
not gate_166(G2511,G2505);
not gate_167(G2512,G2508);
nand gate_168(G2518,G2459,G2460);
buf gate_169(G2551,G1344);
buf gate_170(G2559,G1351);
buf gate_171(G2567,G1959);
buf gate_172(G2575,G1964);
buf gate_173(G2583,G1969);
buf gate_174(G2591,G1974);
buf gate_175(G2599,G1979);
buf gate_176(G2607,G1984);
buf gate_177(G2615,G1989);
buf gate_178(G2623,G1994);
not gate_179(G2705,G2699);
not gate_180(G2706,G2702);
buf gate_181(G2735,G1999);
buf gate_182(G2743,G2070);
buf gate_183(G2751,G2076);
buf gate_184(G2759,G2082);
buf gate_185(G2767,G2088);
buf gate_186(G2775,G2094);
not gate_187(G217,G216);
and gate_188(G550,G2106,G1253);
and gate_189(G552,G567,G1256);
buf gate_190(G325,G558);
or gate_191(G894,G881,G882);
nand gate_192(G1498,G2474,G2477);
nand gate_193(G1507,G2482,G2485);
nand gate_194(G1508,G2479,G2486);
nand gate_195(G1516,G2490,G2493);
nand gate_196(G1517,G2487,G2494);
nand gate_197(G1775,G2678,G2681);
nand gate_198(G1784,G2686,G2689);
nand gate_199(G1785,G2683,G2690);
nand gate_200(G1793,G2694,G2697);
nand gate_201(G1794,G2691,G2698);
nand gate_202(G2469,G2464,G2467);
nand gate_203(G2470,G2461,G2468);
nand gate_204(G2503,G2498,G2501);
nand gate_205(G2504,G2495,G2502);
nand gate_206(G2513,G2508,G2511);
nand gate_207(G2514,G2505,G2512);
nand gate_208(G2707,G2702,G2705);
nand gate_209(G2708,G2699,G2706);
not gate_210(G261,G558);
not gate_211(G551,G550);
not gate_212(G553,G552);
and gate_213(G818,G93,G784,G807);
and gate_214(G819,G55,G772,G807);
and gate_215(G820,G67,G784,G795);
and gate_216(G822,G81,G784,G807);
and gate_217(G823,G43,G772,G807);
and gate_218(G824,G56,G784,G795);
and gate_219(G826,G92,G784,G807);
and gate_220(G827,G54,G772,G807);
and gate_221(G828,G66,G784,G795);
and gate_222(G830,G91,G784,G807);
and gate_223(G831,G53,G772,G807);
and gate_224(G832,G65,G784,G795);
and gate_225(G834,G90,G784,G807);
and gate_226(G835,G52,G772,G807);
and gate_227(G836,G64,G784,G795);
and gate_228(G1307,G89,G1273,G1296);
and gate_229(G1308,G51,G1261,G1296);
and gate_230(G1309,G63,G1273,G1284);
and gate_231(G1311,G88,G1273,G1296);
and gate_232(G1312,G50,G1261,G1296);
and gate_233(G1313,G62,G1273,G1284);
and gate_234(G1315,G87,G1273,G1296);
and gate_235(G1316,G49,G1261,G1296);
and gate_236(G1317,G1273,G1284);
and gate_237(G1319,G86,G1273,G1296);
and gate_238(G1320,G48,G1261,G1296);
and gate_239(G1321,G61,G1273,G1284);
and gate_240(G1323,G85,G1273,G1296);
and gate_241(G1324,G47,G1261,G1296);
and gate_242(G1325,G60,G1273,G1284);
and gate_243(G1441,G138,G1406,G1430);
and gate_244(G1442,G102,G1394,G1430);
and gate_245(G1443,G126,G1406,G1418);
and gate_246(G1445,G137,G1406,G1430);
and gate_247(G1446,G101,G1394,G1430);
and gate_248(G1447,G125,G1406,G1418);
and gate_249(G1449,G136,G1406,G1430);
and gate_250(G1450,G100,G1394,G1430);
and gate_251(G1451,G124,G1406,G1418);
and gate_252(G1453,G135,G1406,G1430);
and gate_253(G1454,G99,G1394,G1430);
and gate_254(G1455,G123,G1406,G1418);
and gate_255(G1457,G1406,G1430);
and gate_256(G1458,G1394,G1430);
and gate_257(G1459,G1406,G1418);
not gate_258(G1481,G1477);
not gate_259(G1490,G1486);
nand gate_260(G1500,G1498,G1499);
nand gate_261(G1509,G1507,G1508);
nand gate_262(G1518,G1516,G1517);
buf gate_263(G1521,G1495);
buf gate_264(G1525,G1495);
not gate_265(G2557,G2551);
not gate_266(G2565,G2559);
not gate_267(G2573,G2567);
not gate_268(G2581,G2575);
not gate_269(G2589,G2583);
not gate_270(G2597,G2591);
not gate_271(G2605,G2599);
not gate_272(G2613,G2607);
not gate_273(G2621,G2615);
not gate_274(G2629,G2623);
and gate_275(G1678,G142,G1643,G1667);
and gate_276(G1679,G106,G1631,G1667);
and gate_277(G1680,G130,G1643,G1655);
and gate_278(G1682,G131,G1643,G1667);
and gate_279(G1683,G95,G1631,G1667);
and gate_280(G1684,G119,G1643,G1655);
and gate_281(G1686,G141,G1643,G1667);
and gate_282(G1687,G105,G1631,G1667);
and gate_283(G1688,G129,G1643,G1655);
and gate_284(G1690,G140,G1643,G1667);
and gate_285(G1691,G104,G1631,G1667);
and gate_286(G1692,G128,G1643,G1655);
and gate_287(G1694,G139,G1643,G1667);
and gate_288(G1695,G103,G1631,G1667);
and gate_289(G1696,G127,G1643,G1655);
and gate_290(G1734,G19,G1716);
and gate_291(G1736,G4,G1716);
and gate_292(G1738,G20,G1716);
and gate_293(G1740,G5,G1716);
and gate_294(G1742,G21,G1728);
and gate_295(G1744,G22,G1728);
and gate_296(G1746,G23,G1728);
and gate_297(G1748,G6,G1728);
and gate_298(G1750,G24,G1728);
nand gate_299(G1777,G1775,G1776);
nand gate_300(G1786,G1784,G1785);
nand gate_301(G1795,G1793,G1794);
and gate_302(G2023,G25,G2007);
and gate_303(G2025,G32,G2007);
and gate_304(G2027,G26,G2007);
and gate_305(G2029,G33,G2007);
and gate_306(G2031,G27,G2018);
and gate_307(G2033,G34,G2018);
and gate_308(G2035,G35,G2018);
and gate_309(G2037,G28,G2018);
not gate_310(G2741,G2735);
not gate_311(G2749,G2743);
not gate_312(G2757,G2751);
not gate_313(G2765,G2759);
not gate_314(G2773,G2767);
not gate_315(G2781,G2775);
nand gate_316(G2515,G2469,G2470);
not gate_317(G2522,G2518);
nand gate_318(G2525,G2513,G2514);
nand gate_319(G2528,G2503,G2504);
nand gate_320(G2730,G2707,G2708);
and gate_321(G554,G551,G553);
or gate_322(G838,G818,G819,G820,G821);
or gate_323(G841,G822,G823,G824,G825);
or gate_324(G846,G826,G827,G828,G829);
or gate_325(G854,G830,G831,G832,G833);
or gate_326(G857,G834,G835,G836,G837);
or gate_327(G1327,G1307,G1308,G1309,G1310);
or gate_328(G1329,G1311,G1312,G1313,G1314);
or gate_329(G1331,G1315,G1316,G1317,G1318);
or gate_330(G1333,G1319,G1320,G1321,G1322);
or gate_331(G1335,G1323,G1324,G1325,G1326);
or gate_332(G1461,G1441,G1442,G1443,G1444);
or gate_333(G1464,G1445,G1446,G1447,G1448);
or gate_334(G1467,G1449,G1450,G1451,G1452);
or gate_335(G1470,G1453,G1454,G1455,G1456);
or gate_336(G1473,G1457,G1458,G1459,G1460);
or gate_337(G1698,G1682,G1683,G1684,G1685);
or gate_338(G1701,G1686,G1687,G1688,G1689);
or gate_339(G1704,G1690,G1691,G1692,G1693);
or gate_340(G1707,G1694,G1695,G1696,G1697);
or gate_341(G2634,G1678,G1679,G1680,G1681);
buf gate_342(G319,G554);
not gate_343(G1504,G1500);
not gate_344(G1513,G1509);
not gate_345(G1524,G1521);
not gate_346(G1528,G1525);
buf gate_347(G1529,G1518);
buf gate_348(G1533,G1518);
and gate_349(G1538,G1486,G1477,G1521);
and gate_350(G1541,G1490,G1481,G1525);
not gate_351(G1781,G1777);
not gate_352(G1790,G1786);
buf gate_353(G1806,G1795);
buf gate_354(G1810,G1795);
not gate_355(G2734,G2730);
not gate_356(G2521,G2515);
nand gate_357(G2524,G2515,G2522);
not gate_358(G2531,G2525);
not gate_359(G2532,G2528);
and gate_360(G144,G838,G860);
and gate_361(G147,G846,G860);
and gate_362(G152,G841,G860);
not gate_363(G160,G1464);
not gate_364(G162,G1467);
not gate_365(G164,G1461);
not gate_366(G166,G1329);
not gate_367(G168,G1327);
not gate_368(G171,G857);
and gate_369(G175,G480,G483,G36,G554);
and gate_370(G187,G480,G483,G554,G547);
buf gate_371(G516,G838);
not gate_372(G852,G846);
and gate_373(G885,G841,G875);
and gate_374(G887,G846,G875);
and gate_375(G893,G1327,G868);
not gate_376(G1028,G838);
not gate_377(G1031,G841);
not gate_378(G1035,G846);
buf gate_379(G1041,G854);
buf gate_380(G1049,G857);
buf gate_381(G1057,G1327);
buf gate_382(G1060,G1329);
buf gate_383(G1066,G1331);
buf gate_384(G1072,G1333);
buf gate_385(G1078,G1335);
nand gate_386(G1213,G2099,G1470);
nand gate_387(G1218,G2103,G1473);
buf gate_388(G1250,G1704);
and gate_389(G1387,G1461,G1385);
not gate_390(G1389,G1464);
and gate_391(G1537,G1481,G1486,G1524);
and gate_392(G1540,G1477,G1490,G1528);
and gate_393(G1735,G841,G1710);
and gate_394(G1737,G846,G1710);
and gate_395(G1739,G854,G1710);
and gate_396(G1741,G857,G1710);
and gate_397(G1743,G1327,G1721);
and gate_398(G1745,G1329,G1721);
and gate_399(G1747,G1331,G1721);
and gate_400(G1749,G1333,G1721);
and gate_401(G1751,G1335,G1721);
not gate_402(G2638,G2634);
and gate_403(G2024,G1698,G2001);
and gate_404(G2026,G1701,G2001);
and gate_405(G2028,G1704,G2001);
and gate_406(G2030,G1707,G2001);
and gate_407(G2032,G1461,G2012);
and gate_408(G2034,G1464,G2012);
and gate_409(G2036,G1467,G2012);
and gate_410(G2038,G1470,G2012);
buf gate_411(G2154,G841);
nand gate_412(G2523,G2518,G2521);
nand gate_413(G2533,G2528,G2531);
nand gate_414(G2534,G2525,G2532);
buf gate_415(G2631,G1698);
buf gate_416(G2639,G1704);
buf gate_417(G2642,G1701);
buf gate_418(G2647,G1461);
buf gate_419(G2650,G1707);
buf gate_420(G2655,G1467);
buf gate_421(G2658,G1464);
buf gate_422(G2665,G1473);
buf gate_423(G2668,G1470);
or gate_424(G153,G865,G152);
not gate_425(G176,G175);
not gate_426(G188,G187);
buf gate_427(G299,G1041);
buf gate_428(G301,G1049);
buf gate_429(G286,G1057);
buf gate_430(G303,G1060);
buf gate_431(G288,G1066);
buf gate_432(G305,G1072);
buf gate_433(G290,G1078);
not gate_434(G1532,G1529);
not gate_435(G1536,G1533);
nor gate_436(G1539,G1537,G1538);
nor gate_437(G1542,G1540,G1541);
and gate_438(G1544,G1509,G1500,G1529);
and gate_439(G1547,G1513,G1504,G1533);
or gate_440(G2065,G2037,G2038);
not gate_441(G1809,G1806);
not gate_442(G1813,G1810);
and gate_443(G1821,G1786,G1777,G1806);
and gate_444(G1824,G1790,G1781,G1810);
nand gate_445(G2538,G2523,G2524);
nand gate_446(G2546,G2533,G2534);
or gate_447(G2554,G1734,G1735);
or gate_448(G2562,G1736,G1737);
or gate_449(G2570,G1738,G1739);
or gate_450(G2578,G1740,G1741);
or gate_451(G2586,G1742,G1743);
or gate_452(G2594,G1744,G1745);
or gate_453(G2602,G1746,G1747);
or gate_454(G2610,G1748,G1749);
or gate_455(G2618,G1750,G1751);
or gate_456(G2626,G2023,G2024);
or gate_457(G2738,G2025,G2026);
or gate_458(G2746,G2027,G2028);
or gate_459(G2754,G2029,G2030);
or gate_460(G2762,G2031,G2032);
or gate_461(G2770,G2033,G2034);
or gate_462(G2778,G2035,G2036);
and gate_463(G456,G1389,G1387,G40);
not gate_464(G466,G1387);
nand gate_465(G562,G560,G852);
and gate_466(G883,G516,G875);
and gate_467(G889,G1049,G868);
and gate_468(G891,G1041,G875);
not gate_469(G1043,G1041);
not gate_470(G1051,G1049);
not gate_471(G1062,G1060);
not gate_472(G1068,G1066);
not gate_473(G1074,G1072);
not gate_474(G1080,G1078);
and gate_475(G1225,G2099,G1213);
and gate_476(G1227,G1213,G1470);
and gate_477(G1232,G2103,G1218);
and gate_478(G1234,G1218,G1473);
and gate_479(G1543,G1504,G1509,G1532);
and gate_480(G1546,G1500,G1513,G1536);
not gate_481(G2637,G2631);
nand gate_482(G1753,G2631,G2638);
not gate_483(G2645,G2639);
not gate_484(G2646,G2642);
not gate_485(G2653,G2647);
not gate_486(G2654,G2650);
and gate_487(G1820,G1781,G1786,G1809);
and gate_488(G1823,G1777,G1790,G1813);
buf gate_489(G2107,G1031);
buf gate_490(G2110,G1028);
buf gate_491(G2118,G1035);
not gate_492(G2123,G1057);
not gate_493(G2151,G852);
not gate_494(G2158,G2154);
buf gate_495(G2161,G1031);
buf gate_496(G2164,G1028);
buf gate_497(G2172,G1035);
buf gate_498(G2235,G516);
buf gate_499(G2262,G1035);
buf gate_500(G2350,G1035);
nand gate_501(G2535,G1542,G1539);
not gate_502(G2661,G2655);
not gate_503(G2662,G2658);
not gate_504(G2671,G2665);
not gate_505(G2672,G2668);
and gate_506(G468,G40,G1389,G466);
or gate_507(G897,G887,G889);
or gate_508(G898,G891,G893);
or gate_509(G1228,G1225,G1227);
or gate_510(G1235,G1232,G1234);
nor gate_511(G1545,G1543,G1544);
nor gate_512(G1548,G1546,G1547);
not gate_513(G2542,G2538);
not gate_514(G2550,G2546);
nand gate_515(G1561,G2554,G2557);
not gate_516(G2558,G2554);
nand gate_517(G1565,G2562,G2565);
not gate_518(G2566,G2562);
nand gate_519(G1569,G2570,G2573);
not gate_520(G2574,G2570);
nand gate_521(G1573,G2578,G2581);
not gate_522(G2582,G2578);
nand gate_523(G1577,G2586,G2589);
not gate_524(G2590,G2586);
nand gate_525(G1581,G2594,G2597);
not gate_526(G2598,G2594);
nand gate_527(G1585,G2602,G2605);
not gate_528(G2606,G2602);
nand gate_529(G1589,G2610,G2613);
not gate_530(G2614,G2610);
nand gate_531(G1593,G2618,G2621);
not gate_532(G2622,G2618);
nand gate_533(G1597,G2626,G2629);
not gate_534(G2630,G2626);
nand gate_535(G1752,G2634,G2637);
nand gate_536(G1761,G2642,G2645);
nand gate_537(G1762,G2639,G2646);
nand gate_538(G1770,G2650,G2653);
nand gate_539(G1771,G2647,G2654);
nor gate_540(G1822,G1820,G1821);
nor gate_541(G1825,G1823,G1824);
nand gate_542(G2039,G2738,G2741);
not gate_543(G2742,G2738);
nand gate_544(G2043,G2746,G2749);
not gate_545(G2750,G2746);
nand gate_546(G2047,G2754,G2757);
not gate_547(G2758,G2754);
nand gate_548(G2051,G2762,G2765);
not gate_549(G2766,G2762);
nand gate_550(G2055,G2770,G2773);
not gate_551(G2774,G2770);
nand gate_552(G2059,G2778,G2781);
not gate_553(G2782,G2778);
nand gate_554(G2663,G2658,G2661);
nand gate_555(G2664,G2655,G2662);
nand gate_556(G2673,G2668,G2671);
nand gate_557(G2674,G2665,G2672);
and gate_558(G146,G562,G865);
not gate_559(G462,G456);
not gate_560(G2113,G2107);
not gate_561(G2114,G2110);
not gate_562(G2122,G2118);
not gate_563(G2129,G2123);
buf gate_564(G592,G562);
not gate_565(G2167,G2161);
not gate_566(G2168,G2164);
not gate_567(G2176,G2172);
not gate_568(G2241,G2235);
not gate_569(G2266,G2262);
not gate_570(G743,G456);
buf gate_571(G749,G456);
and gate_572(G886,G562,G868);
buf gate_573(G284,G897);
buf gate_574(G321,G897);
buf gate_575(G297,G898);
buf gate_576(G280,G898);
buf gate_577(G995,G456);
not gate_578(G1006,G456);
nand gate_579(G1550,G2535,G2542);
not gate_580(G2354,G2350);
not gate_581(G2541,G2535);
nand gate_582(G1562,G2551,G2558);
nand gate_583(G1566,G2559,G2566);
nand gate_584(G1570,G2567,G2574);
nand gate_585(G1574,G2575,G2582);
nand gate_586(G1578,G2583,G2590);
nand gate_587(G1582,G2591,G2598);
nand gate_588(G1586,G2599,G2606);
nand gate_589(G1590,G2607,G2614);
nand gate_590(G1594,G2615,G2622);
nand gate_591(G1598,G2623,G2630);
nand gate_592(G1754,G1752,G1753);
nand gate_593(G1763,G1761,G1762);
nand gate_594(G1772,G1770,G1771);
nand gate_595(G2040,G2735,G2742);
nand gate_596(G2044,G2743,G2750);
nand gate_597(G2048,G2751,G2758);
nand gate_598(G2052,G2759,G2766);
nand gate_599(G2056,G2767,G2774);
nand gate_600(G2060,G2775,G2782);
buf gate_601(G2115,G1043);
buf gate_602(G2126,G1051);
buf gate_603(G2131,G1068);
buf gate_604(G2134,G1062);
buf gate_605(G2141,G1080);
buf gate_606(G2144,G1074);
not gate_607(G2157,G2151);
nand gate_608(G2160,G2151,G2158);
buf gate_609(G2169,G1043);
buf gate_610(G2177,G1068);
buf gate_611(G2180,G1062);
buf gate_612(G2187,G1080);
buf gate_613(G2190,G1074);
not gate_614(G2207,G562);
buf gate_615(G2254,G1043);
buf gate_616(G2334,G1051);
buf gate_617(G2342,G1043);
buf gate_618(G2422,G1051);
nand gate_619(G2543,G1548,G1545);
nand gate_620(G2709,G2673,G2674);
nand gate_621(G2712,G2663,G2664);
nand gate_622(G2727,G1825,G1822);
or gate_623(G148,G146,G147);
nand gate_624(G569,G2110,G2113);
nand gate_625(G570,G2107,G2114);
nand gate_626(G599,G2164,G2167);
nand gate_627(G600,G2161,G2168);
or gate_628(G896,G885,G886);
nand gate_629(G1549,G2538,G2541);
not gate_630(G1243,G1228);
not gate_631(G1245,G1235);
buf gate_632(G1257,G468);
buf gate_633(G1258,G468);
nand gate_634(G1563,G1561,G1562);
nand gate_635(G1567,G1565,G1566);
nand gate_636(G1571,G1569,G1570);
nand gate_637(G1575,G1573,G1574);
nand gate_638(G1579,G1577,G1578);
nand gate_639(G1583,G1581,G1582);
nand gate_640(G1587,G1585,G1586);
nand gate_641(G1591,G1589,G1590);
nand gate_642(G1595,G1593,G1594);
nand gate_643(G1599,G1597,G1598);
nand gate_644(G2041,G2039,G2040);
nand gate_645(G2045,G2043,G2044);
nand gate_646(G2049,G2047,G2048);
nand gate_647(G2053,G2051,G2052);
nand gate_648(G2057,G2055,G2056);
nand gate_649(G2061,G2059,G2060);
nand gate_650(G2159,G2154,G2157);
buf gate_651(G475,G462);
and gate_652(G490,G1078,G743);
and gate_653(G496,G1698,G743);
and gate_654(G502,G1701,G743);
and gate_655(G508,G1250,G743);
and gate_656(G765,G1057,G749);
and gate_657(G769,G1060,G749);
nand gate_658(G571,G569,G570);
not gate_659(G2121,G2115);
nand gate_660(G579,G2115,G2122);
nand gate_661(G587,G2126,G2129);
not gate_662(G2130,G2126);
not gate_663(G596,G592);
nand gate_664(G601,G599,G600);
not gate_665(G2175,G2169);
nand gate_666(G609,G2169,G2176);
not gate_667(G2258,G2254);
and gate_668(G1014,G1057,G995);
and gate_669(G1018,G1060,G995);
and gate_670(G717,G1078,G1006);
and gate_671(G723,G1698,G1006);
and gate_672(G729,G1701,G1006);
and gate_673(G735,G1250,G1006);
not gate_674(G753,G749);
buf gate_675(G282,G896);
buf gate_676(G323,G896);
not gate_677(G2338,G2334);
not gate_678(G999,G995);
nand gate_679(G1091,G1549,G1550);
not gate_680(G2346,G2342);
not gate_681(G2426,G2422);
buf gate_682(G1337,G462);
not gate_683(G2549,G2543);
nand gate_684(G1552,G2543,G2550);
not gate_685(G1600,G1599);
not gate_686(G1596,G1595);
not gate_687(G1592,G1591);
not gate_688(G1588,G1587);
not gate_689(G1584,G1583);
not gate_690(G1580,G1579);
not gate_691(G1576,G1575);
not gate_692(G1572,G1571);
not gate_693(G1568,G1567);
not gate_694(G1564,G1563);
not gate_695(G2062,G2061);
not gate_696(G2058,G2057);
not gate_697(G2054,G2053);
not gate_698(G2050,G2049);
not gate_699(G2046,G2045);
not gate_700(G2042,G2041);
not gate_701(G1758,G1754);
not gate_702(G1767,G1763);
buf gate_703(G1798,G1772);
buf gate_704(G1802,G1772);
not gate_705(G2733,G2727);
nand gate_706(G1829,G2727,G2734);
not gate_707(G2137,G2131);
not gate_708(G2138,G2134);
not gate_709(G2147,G2141);
not gate_710(G2148,G2144);
not gate_711(G2183,G2177);
not gate_712(G2184,G2180);
not gate_713(G2193,G2187);
not gate_714(G2194,G2190);
nand gate_715(G2210,G2159,G2160);
not gate_716(G2213,G2207);
not gate_717(G2715,G2709);
not gate_718(G2716,G2712);
and gate_719(G1094,G1235,G1245);
and gate_720(G1096,G1228,G1243);
nand gate_721(G578,G2118,G2121);
nand gate_722(G588,G2123,G2130);
nand gate_723(G608,G2172,G2175);
buf gate_724(G742,G1257);
buf gate_725(G1005,G1257);
not gate_726(G1092,G1091);
nand gate_727(G1551,G2546,G2549);
and gate_728(G1554,G1600,G1596,G1592,G1588,G1584);
and gate_729(G1555,G1580,G1576,G1572,G1568,G1564);
and gate_730(G1557,G2065,G2062);
and gate_731(G1558,G2058,G2054,G2050,G2046,G2042);
nand gate_732(G1828,G2730,G2733);
buf gate_733(G1845,G1258);
buf gate_734(G1907,G1258);
nand gate_735(G2139,G2134,G2137);
nand gate_736(G2140,G2131,G2138);
nand gate_737(G2149,G2144,G2147);
nand gate_738(G2150,G2141,G2148);
nand gate_739(G2185,G2180,G2183);
nand gate_740(G2186,G2177,G2184);
nand gate_741(G2195,G2190,G2193);
nand gate_742(G2196,G2187,G2194);
nand gate_743(G2717,G2712,G2715);
nand gate_744(G2718,G2709,G2716);
or gate_745(G154,G1094,G1245);
or gate_746(G155,G1096,G1243);
and gate_747(G763,G1057,G753);
and gate_748(G767,G1060,G753);
and gate_749(G531,G1066,G753);
and gate_750(G537,G1072,G753);
not gate_751(G575,G571);
nand gate_752(G580,G578,G579);
nand gate_753(G589,G587,G588);
not gate_754(G605,G601);
nand gate_755(G610,G608,G609);
and gate_756(G1012,G1057,G999);
and gate_757(G1016,G1060,G999);
and gate_758(G705,G1066,G999);
and gate_759(G711,G1072,G999);
and gate_760(G1093,G1092,G14);
buf gate_761(G1355,G475);
nand gate_762(G1553,G1551,G1552);
and gate_763(G1556,G1554,G1555);
and gate_764(G1559,G1557,G1558);
buf gate_765(G1601,G1337);
not gate_766(G1801,G1798);
not gate_767(G1805,G1802);
and gate_768(G1815,G1763,G1754,G1798);
and gate_769(G1818,G1767,G1758,G1802);
nand gate_770(G1830,G1828,G1829);
buf gate_771(G1836,G475);
buf gate_772(G1850,G475);
buf gate_773(G1898,G1337);
buf gate_774(G1912,G1337);
nand gate_775(G2197,G2149,G2150);
nand gate_776(G2200,G2139,G2140);
not gate_777(G2214,G2210);
nand gate_778(G2215,G2210,G2213);
nand gate_779(G2217,G2195,G2196);
nand gate_780(G2220,G2185,G2186);
nand gate_781(G2722,G2717,G2718);
nand gate_782(G156,G154,G155);
and gate_783(G492,G490,G742);
and gate_784(G498,G496,G742);
and gate_785(G504,G502,G742);
and gate_786(G510,G508,G742);
or gate_787(G519,G763,G765);
or gate_788(G525,G767,G769);
and gate_789(G533,G531,G748);
and gate_790(G539,G537,G748);
or gate_791(G693,G1012,G1014);
or gate_792(G699,G1016,G1018);
and gate_793(G707,G705,G994);
and gate_794(G713,G711,G994);
and gate_795(G719,G717,G1005);
and gate_796(G725,G723,G1005);
and gate_797(G731,G729,G1005);
and gate_798(G737,G735,G1005);
buf gate_799(G401,G1093);
and gate_800(G1560,G1556,G1559,G894);
and gate_801(G1814,G1758,G1763,G1801);
and gate_802(G1817,G1754,G1767,G1805);
nand gate_803(G2216,G2207,G2214);
not gate_804(G227,G1830);
not gate_805(G229,G1553);
not gate_806(G493,G492);
not gate_807(G499,G498);
not gate_808(G505,G504);
not gate_809(G511,G510);
and gate_810(G521,G519,G748);
and gate_811(G527,G525,G748);
not gate_812(G534,G533);
not gate_813(G540,G539);
not gate_814(G584,G580);
buf gate_815(G613,G589);
buf gate_816(G617,G589);
buf gate_817(G621,G610);
buf gate_818(G625,G610);
and gate_819(G676,G1344,G1355);
and gate_820(G695,G693,G994);
and gate_821(G701,G699,G994);
not gate_822(G708,G707);
not gate_823(G714,G713);
not gate_824(G720,G719);
not gate_825(G726,G725);
not gate_826(G732,G731);
not gate_827(G738,G737);
not gate_828(G1087,G1093);
and gate_829(G1108,G1344,G1601);
not gate_830(G1361,G1355);
and gate_831(G1369,G1351,G1355);
and gate_832(G1373,G1959,G1355);
and gate_833(G1377,G1964,G1355);
buf gate_834(G311,G1560);
not gate_835(G1607,G1601);
and gate_836(G1615,G1351,G1601);
and gate_837(G1619,G1959,G1601);
and gate_838(G1623,G1964,G1601);
nor gate_839(G1816,G1814,G1815);
nor gate_840(G1819,G1817,G1818);
not gate_841(G2726,G2722);
not gate_842(G1842,G1836);
and gate_843(G1858,G1969,G1836);
and gate_844(G1863,G1974,G1836);
and gate_845(G1866,G1979,G1836);
and gate_846(G1868,G1984,G1836);
and gate_847(G1870,G1989,G1850);
and gate_848(G1872,G1994,G1850);
and gate_849(G1874,G1999,G1850);
and gate_850(G1876,G2070,G1850);
not gate_851(G1904,G1898);
and gate_852(G1920,G1969,G1898);
and gate_853(G1925,G1974,G1898);
and gate_854(G1928,G1979,G1898);
and gate_855(G1930,G1984,G1898);
and gate_856(G1932,G1989,G1912);
and gate_857(G1934,G1994,G1912);
and gate_858(G1936,G1999,G1912);
and gate_859(G1938,G2070,G1912);
not gate_860(G2203,G2197);
not gate_861(G2204,G2200);
not gate_862(G2223,G2217);
not gate_863(G2224,G2220);
nand gate_864(G2238,G2215,G2216);
not gate_865(G150,G1560);
not gate_866(G522,G521);
not gate_867(G528,G527);
not gate_868(G696,G695);
not gate_869(G702,G701);
and gate_870(G1881,G1866,G1831);
and gate_871(G1883,G1868,G1831);
and gate_872(G1885,G1870,G1845);
and gate_873(G1887,G1872,G1845);
and gate_874(G1889,G1874,G1845);
and gate_875(G1891,G1876,G1845);
and gate_876(G1943,G1928,G1893);
and gate_877(G1945,G1930,G1893);
and gate_878(G1947,G1932,G1907);
and gate_879(G1949,G1934,G1907);
and gate_880(G1951,G1936,G1907);
and gate_881(G1953,G1938,G1907);
nand gate_882(G2205,G2200,G2203);
nand gate_883(G2206,G2197,G2204);
nand gate_884(G2225,G2220,G2223);
nand gate_885(G2226,G2217,G2224);
nand gate_886(G2719,G1819,G1816);
not gate_887(G616,G613);
not gate_888(G620,G617);
not gate_889(G624,G621);
not gate_890(G628,G625);
and gate_891(G630,G580,G571,G613);
and gate_892(G633,G584,G575,G617);
and gate_893(G636,G601,G592,G621);
and gate_894(G639,G605,G596,G625);
nand gate_895(G645,G2238,G2241);
not gate_896(G2242,G2238);
and gate_897(G675,G1999,G1361);
and gate_898(G1107,G1999,G1607);
and gate_899(G1368,G2070,G1361);
and gate_900(G1371,G2076,G1361);
and gate_901(G1375,G2082,G1361);
and gate_902(G1614,G2070,G1607);
and gate_903(G1617,G2076,G1607);
and gate_904(G1621,G2082,G1607);
and gate_905(G1856,G2088,G1842);
and gate_906(G1861,G2094,G1842);
and gate_907(G1918,G2088,G1904);
and gate_908(G1923,G2094,G1904);
nand gate_909(G2230,G2205,G2206);
nand gate_910(G2246,G2225,G2226);
buf gate_911(G2270,G511);
buf gate_912(G2278,G505);
buf gate_913(G2286,G499);
buf gate_914(G2294,G493);
buf gate_915(G2302,G540);
buf gate_916(G2310,G534);
buf gate_917(G2358,G738);
buf gate_918(G2366,G732);
buf gate_919(G2374,G726);
buf gate_920(G2382,G720);
buf gate_921(G2390,G714);
buf gate_922(G2398,G708);
and gate_923(G629,G575,G580,G616);
and gate_924(G632,G571,G584,G620);
and gate_925(G635,G596,G601,G624);
and gate_926(G638,G592,G605,G628);
nand gate_927(G646,G2235,G2242);
or gate_928(G677,G675,G676);
nand gate_929(G1827,G2719,G2726);
and gate_930(G907,G1891,G511);
and gate_931(G915,G1889,G505);
and gate_932(G922,G1887,G499);
and gate_933(G924,G493,G1885);
and gate_934(G937,G1883,G540);
and gate_935(G946,G1881,G534);
or gate_936(G1109,G1107,G1108);
and gate_937(G1125,G1953,G738);
and gate_938(G1133,G1951,G732);
and gate_939(G1140,G1949,G726);
and gate_940(G1142,G720,G1947);
and gate_941(G1155,G1945,G714);
and gate_942(G1164,G1943,G708);
or gate_943(G1378,G1368,G1369);
or gate_944(G1380,G1371,G1373);
or gate_945(G1382,G1375,G1377);
or gate_946(G1624,G1614,G1615);
or gate_947(G1626,G1617,G1619);
or gate_948(G1628,G1621,G1623);
not gate_949(G2725,G2719);
or gate_950(G1859,G1856,G1858);
or gate_951(G1864,G1861,G1863);
or gate_952(G1921,G1918,G1920);
or gate_953(G1926,G1923,G1925);
buf gate_954(G2267,G1891);
buf gate_955(G2275,G1889);
buf gate_956(G2283,G1887);
buf gate_957(G2291,G1885);
buf gate_958(G2299,G1883);
buf gate_959(G2307,G1881);
buf gate_960(G2318,G528);
buf gate_961(G2326,G522);
buf gate_962(G2355,G1953);
buf gate_963(G2363,G1951);
buf gate_964(G2371,G1949);
buf gate_965(G2379,G1947);
buf gate_966(G2387,G1945);
buf gate_967(G2395,G1943);
buf gate_968(G2406,G702);
buf gate_969(G2414,G696);
nand gate_970(G647,G645,G646);
nor gate_971(G631,G629,G630);
nor gate_972(G634,G632,G633);
nor gate_973(G637,G635,G636);
nor gate_974(G640,G638,G639);
not gate_975(G2234,G2230);
not gate_976(G2250,G2246);
and gate_977(G679,G677,G1031);
nand gate_978(G1826,G2722,G2725);
not gate_979(G2274,G2270);
not gate_980(G2282,G2278);
not gate_981(G2290,G2286);
not gate_982(G2298,G2294);
not gate_983(G2306,G2302);
not gate_984(G2314,G2310);
and gate_985(G1110,G1109,G1031);
not gate_986(G2362,G2358);
not gate_987(G2370,G2366);
not gate_988(G2378,G2374);
not gate_989(G2386,G2382);
not gate_990(G2394,G2390);
not gate_991(G2402,G2398);
and gate_992(G1877,G1859,G1831);
and gate_993(G1879,G1864,G1831);
and gate_994(G1939,G1921,G1893);
and gate_995(G1941,G1926,G1893);
and gate_996(G143,G647,G865);
and gate_997(G671,G1380,G1043);
and gate_998(G674,G1378,G1035);
nand gate_999(G686,G1826,G1827);
not gate_1000(G2273,G2267);
nand gate_1001(G900,G2267,G2274);
not gate_1002(G2281,G2275);
nand gate_1003(G909,G2275,G2282);
not gate_1004(G2289,G2283);
nand gate_1005(G917,G2283,G2290);
not gate_1006(G2297,G2291);
nand gate_1007(G926,G2291,G2298);
not gate_1008(G2305,G2299);
nand gate_1009(G929,G2299,G2306);
not gate_1010(G2313,G2307);
nand gate_1011(G939,G2307,G2314);
not gate_1012(G2322,G2318);
not gate_1013(G2330,G2326);
and gate_1014(G967,G1382,G1051);
and gate_1015(G1104,G1626,G1043);
and gate_1016(G1106,G1624,G1035);
not gate_1017(G2361,G2355);
nand gate_1018(G1118,G2355,G2362);
not gate_1019(G2369,G2363);
nand gate_1020(G1127,G2363,G2370);
not gate_1021(G2377,G2371);
nand gate_1022(G1135,G2371,G2378);
not gate_1023(G2385,G2379);
nand gate_1024(G1144,G2379,G2386);
not gate_1025(G2393,G2387);
nand gate_1026(G1147,G2387,G2394);
not gate_1027(G2401,G2395);
nand gate_1028(G1157,G2395,G2402);
not gate_1029(G2410,G2406);
not gate_1030(G2418,G2414);
and gate_1031(G1184,G1628,G1051);
nand gate_1032(G2227,G634,G631);
nand gate_1033(G2243,G640,G637);
buf gate_1034(G2251,G1380);
buf gate_1035(G2259,G1378);
buf gate_1036(G2331,G1382);
buf gate_1037(G2339,G1626);
buf gate_1038(G2347,G1624);
buf gate_1039(G2419,G1628);
or gate_1040(G145,G143,G144);
not gate_1041(G687,G686);
nand gate_1042(G899,G2270,G2273);
nand gate_1043(G908,G2278,G2281);
nand gate_1044(G916,G2286,G2289);
nand gate_1045(G925,G2294,G2297);
nand gate_1046(G928,G2302,G2305);
nand gate_1047(G938,G2310,G2313);
and gate_1048(G954,G1879,G528);
and gate_1049(G961,G1877,G522);
nand gate_1050(G1117,G2358,G2361);
nand gate_1051(G1126,G2366,G2369);
nand gate_1052(G1134,G2374,G2377);
nand gate_1053(G1143,G2382,G2385);
nand gate_1054(G1146,G2390,G2393);
nand gate_1055(G1156,G2398,G2401);
and gate_1056(G1172,G1941,G702);
and gate_1057(G1179,G1939,G696);
buf gate_1058(G2315,G1879);
buf gate_1059(G2323,G1877);
buf gate_1060(G2403,G1941);
buf gate_1061(G2411,G1939);
not gate_1062(G2233,G2227);
nand gate_1063(G642,G2227,G2234);
not gate_1064(G2249,G2243);
nand gate_1065(G649,G2243,G2250);
not gate_1066(G2257,G2251);
nand gate_1067(G665,G2251,G2258);
nand gate_1068(G684,G2259,G2266);
not gate_1069(G2265,G2259);
and gate_1070(G688,G687,G487);
nand gate_1071(G901,G899,G900);
nand gate_1072(G910,G908,G909);
nand gate_1073(G918,G916,G917);
nand gate_1074(G927,G925,G926);
nand gate_1075(G930,G928,G929);
nand gate_1076(G940,G938,G939);
not gate_1077(G2337,G2331);
nand gate_1078(G963,G2331,G2338);
not gate_1079(G2345,G2339);
nand gate_1080(G1099,G2339,G2346);
nand gate_1081(G1115,G2347,G2354);
not gate_1082(G2353,G2347);
nand gate_1083(G1119,G1117,G1118);
nand gate_1084(G1128,G1126,G1127);
nand gate_1085(G1136,G1134,G1135);
nand gate_1086(G1145,G1143,G1144);
nand gate_1087(G1148,G1146,G1147);
nand gate_1088(G1158,G1156,G1157);
not gate_1089(G2425,G2419);
nand gate_1090(G1181,G2419,G2426);
nand gate_1091(G641,G2230,G2233);
nand gate_1092(G648,G2246,G2249);
nand gate_1093(G664,G2254,G2257);
nand gate_1094(G683,G2262,G2265);
buf gate_1095(G395,G688);
not gate_1096(G2321,G2315);
nand gate_1097(G948,G2315,G2322);
not gate_1098(G2329,G2323);
nand gate_1099(G956,G2323,G2330);
nand gate_1100(G962,G2334,G2337);
nand gate_1101(G1098,G2342,G2345);
nand gate_1102(G1114,G2350,G2353);
not gate_1103(G2409,G2403);
nand gate_1104(G1166,G2403,G2410);
not gate_1105(G2417,G2411);
nand gate_1106(G1174,G2411,G2418);
nand gate_1107(G1180,G2422,G2425);
nand gate_1108(G643,G641,G642);
nand gate_1109(G650,G648,G649);
nand gate_1110(G666,G664,G665);
nand gate_1111(G681,G683,G684);
not gate_1112(G690,G688);
nand gate_1113(G947,G2318,G2321);
nand gate_1114(G955,G2326,G2329);
nand gate_1115(G964,G962,G963);
and gate_1116(G968,G910,G927,G918,G901);
and gate_1117(G970,G901,G915);
and gate_1118(G971,G910,G901,G922);
and gate_1119(G972,G918,G901,G924,G910);
and gate_1120(G978,G930,G946);
and gate_1121(G979,G940,G930,G954);
nand gate_1122(G1100,G1098,G1099);
nand gate_1123(G1112,G1114,G1115);
nand gate_1124(G1165,G2406,G2409);
nand gate_1125(G1173,G2414,G2417);
nand gate_1126(G1182,G1180,G1181);
and gate_1127(G1185,G1128,G1145,G1136,G1119);
and gate_1128(G1187,G1119,G1133);
and gate_1129(G1188,G1128,G1119,G1140);
and gate_1130(G1189,G1136,G1119,G1142,G1128);
and gate_1131(G1195,G1148,G1164);
and gate_1132(G1196,G1158,G1148,G1172);
not gate_1133(G644,G643);
and gate_1134(G884,G650,G868);
nand gate_1135(G949,G947,G948);
nand gate_1136(G957,G955,G956);
not gate_1137(G969,G968);
or gate_1138(G973,G907,G970,G971,G972);
nand gate_1139(G1167,G1165,G1166);
nand gate_1140(G1175,G1173,G1174);
not gate_1141(G1186,G1185);
or gate_1142(G1190,G1125,G1187,G1188,G1189);
and gate_1143(G680,G666,G674);
and gate_1144(G682,G681,G666,G679);
or gate_1145(G895,G883,G884);
and gate_1146(G1025,G644,G487);
and gate_1147(G1111,G1100,G1106);
and gate_1148(G1113,G1112,G1100,G1110);
or gate_1149(G685,G671,G680,G682);
buf gate_1150(G295,G895);
buf gate_1151(G331,G895);
not gate_1152(G976,G973);
and gate_1153(G977,G940,G964,G949,G930,G957);
and gate_1154(G980,G949,G930,G961,G940);
and gate_1155(G981,G957,G949,G930,G967,G940);
buf gate_1156(G397,G1025);
or gate_1157(G1116,G1104,G1111,G1113);
not gate_1158(G1193,G1190);
and gate_1159(G1194,G1158,G1182,G1167,G1148,G1175);
and gate_1160(G1197,G1167,G1148,G1179,G1158);
and gate_1161(G1198,G1175,G1167,G1148,G1184,G1158);
or gate_1162(G982,G937,G978,G979,G980,G981);
and gate_1163(G983,G977,G685);
nand gate_1164(G988,G976,G969);
not gate_1165(G1027,G1025);
or gate_1166(G1199,G1155,G1195,G1196,G1197,G1198);
and gate_1167(G1200,G1194,G1116);
nand gate_1168(G1205,G1193,G1186);
or gate_1169(G984,G982,G983);
and gate_1170(G1085,G690,G1027,G1830);
or gate_1171(G1201,G1199,G1200);
not gate_1172(G987,G984);
and gate_1173(G990,G988,G984);
not gate_1174(G1204,G1201);
and gate_1175(G1207,G1205,G1201);
and gate_1176(G989,G973,G987);
and gate_1177(G1206,G1190,G1204);
or gate_1178(G991,G989,G990);
or gate_1179(G1208,G1206,G1207);
buf gate_1180(G329,G1208);
nand gate_1181(G1221,G1208,G991);
and gate_1182(G1238,G1208,G1221);
and gate_1183(G1239,G1221,G991);
or gate_1184(G1240,G1238,G1239);
not gate_1185(G1247,G1240);
and gate_1186(G471,G1240,G1247);
or gate_1187(G473,G471,G1247);
not gate_1188(G231,G473);
and gate_1189(G1088,G1553,G1087,G473);
and gate_1190(G1089,G1085,G1088,G554);
buf gate_1191(G308,G1089);
not gate_1192(G225,G1089);
endmodule
