// Verilog File 
module ex1010 (pi0,pi1,pi2,pi3,pi4,pi5,pi6,pi7,pi8,
pi9,po0,po1,po2,po3,po4,po5,po6,po7,po8,
po9);

input pi0,pi1,pi2,pi3,pi4,pi5,pi6,pi7,pi8,
pi9;

output po0,po1,po2,po3,po4,po5,po6,po7,po8,
po9;

wire n20,n21,n22,n23,n24,n25,n26,n27,n28,
n29,n30,n31,n32,n33,n34,n35,n36,n37,n38,
n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,
n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,
n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,
n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,
n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,
n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,
n99,n100,n101,n102,n103,n104,n105,n106,n107,n108,
n109,n110,n111,n112,n113,n114,n115,n116,n117,n118,
n119,n120,n121,n122,n123,n124,n125,n126,n127,n128,
n129,n130,n131,n132,n133,n134,n135,n136,n137,n138,
n139,n140,n141,n142,n143,n144,n145,n146,n147,n148,
n149,n150,n151,n152,n153,n154,n155,n156,n157,n158,
n159,n160,n161,n162,n163,n164,n165,n166,n167,n168,
n169,n170,n171,n172,n173,n174,n175,n176,n177,n178,
n179,n180,n181,n182,n183,n184,n185,n186,n187,n188,
n189,n190,n191,n192,n193,n194,n195,n196,n197,n198,
n199,n200,n201,n202,n203,n204,n205,n206,n207,n208,
n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,
n219,n220,n221,n222,n223,n224,n225,n226,n227,n228,
n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,
n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,
n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,
n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,
n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,
n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,
n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,
n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,
n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,
n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,
n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,
n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,
n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,
n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,
n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,
n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,
n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,
n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,
n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,
n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,
n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,
n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,
n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,
n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,
n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,
n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,
n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,
n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,
n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,
n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,
n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,
n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,
n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,
n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,
n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,
n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,
n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,
n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,
n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,
n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,
n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,
n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,
n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,
n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,
n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,
n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,
n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,
n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,
n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,
n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,
n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,
n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,
n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,
n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,
n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,
n779,n780,n781,n782,n783,n784,n785,n786,n787,n788,
n789,n790,n791,n792,n793,n794,n795,n796,n797,n798,
n799,n800,n801,n802,n803,n804,n805,n806,n807,n808,
n810,n811,n812,n813,n814,n815,n816,n817,n818,n819,
n820,n821,n822,n823,n824,n825,n826,n827,n828,n829,
n830,n831,n832,n833,n834,n835,n836,n837,n838,n839,
n840,n841,n842,n843,n844,n845,n846,n847,n848,n849,
n850,n851,n852,n853,n854,n855,n856,n857,n858,n859,
n860,n861,n862,n863,n864,n865,n866,n867,n868,n869,
n870,n871,n872,n873,n874,n875,n876,n877,n878,n879,
n880,n881,n882,n883,n884,n885,n886,n887,n888,n889,
n890,n891,n892,n893,n894,n895,n896,n897,n898,n899,
n900,n901,n902,n903,n904,n905,n906,n907,n908,n909,
n910,n911,n912,n913,n914,n915,n916,n917,n918,n919,
n920,n921,n922,n923,n924,n925,n926,n927,n928,n929,
n930,n931,n932,n933,n934,n935,n936,n937,n938,n939,
n940,n941,n942,n943,n944,n945,n946,n947,n948,n949,
n950,n951,n952,n953,n954,n955,n956,n957,n958,n959,
n960,n961,n962,n963,n964,n965,n966,n967,n968,n969,
n970,n971,n972,n973,n974,n975,n976,n977,n978,n979,
n980,n981,n982,n983,n984,n985,n986,n987,n988,n989,
n990,n991,n992,n993,n994,n995,n996,n997,n998,n999,
n1000,n1001,n1002,n1003,n1004,n1005,n1006,n1007,n1008,n1009,
n1010,n1011,n1012,n1013,n1014,n1015,n1016,n1017,n1018,n1019,
n1020,n1021,n1022,n1023,n1024,n1025,n1026,n1027,n1028,n1029,
n1030,n1031,n1032,n1033,n1034,n1035,n1036,n1037,n1038,n1039,
n1040,n1041,n1042,n1043,n1044,n1045,n1046,n1047,n1048,n1049,
n1050,n1051,n1052,n1053,n1054,n1055,n1056,n1057,n1058,n1059,
n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,n1069,
n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,n1079,
n1080,n1081,n1082,n1083,n1084,n1085,n1086,n1087,n1088,n1089,
n1090,n1091,n1092,n1093,n1094,n1095,n1096,n1097,n1098,n1099,
n1100,n1101,n1102,n1103,n1104,n1105,n1106,n1107,n1108,n1109,
n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,n1118,n1119,
n1120,n1121,n1122,n1123,n1124,n1125,n1126,n1127,n1128,n1129,
n1130,n1131,n1132,n1133,n1134,n1135,n1136,n1137,n1138,n1139,
n1140,n1141,n1142,n1143,n1144,n1145,n1146,n1147,n1148,n1149,
n1150,n1151,n1152,n1153,n1154,n1155,n1156,n1157,n1158,n1159,
n1160,n1161,n1162,n1163,n1164,n1165,n1166,n1167,n1168,n1169,
n1170,n1171,n1172,n1173,n1174,n1175,n1176,n1177,n1178,n1179,
n1180,n1181,n1182,n1183,n1184,n1185,n1186,n1187,n1188,n1189,
n1190,n1191,n1192,n1193,n1194,n1195,n1196,n1197,n1198,n1199,
n1200,n1201,n1202,n1203,n1204,n1205,n1206,n1207,n1208,n1209,
n1210,n1211,n1212,n1213,n1214,n1215,n1216,n1217,n1218,n1219,
n1220,n1221,n1222,n1223,n1224,n1225,n1226,n1227,n1228,n1229,
n1230,n1231,n1232,n1233,n1234,n1235,n1236,n1237,n1238,n1239,
n1240,n1241,n1242,n1243,n1244,n1245,n1246,n1247,n1248,n1249,
n1250,n1251,n1252,n1253,n1254,n1255,n1256,n1257,n1258,n1259,
n1260,n1261,n1262,n1263,n1264,n1265,n1266,n1267,n1268,n1269,
n1270,n1271,n1272,n1273,n1274,n1275,n1276,n1277,n1278,n1279,
n1280,n1281,n1282,n1283,n1284,n1285,n1286,n1287,n1288,n1289,
n1290,n1291,n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,
n1300,n1301,n1302,n1303,n1304,n1305,n1306,n1307,n1308,n1309,
n1310,n1311,n1312,n1313,n1314,n1315,n1316,n1317,n1318,n1319,
n1320,n1321,n1322,n1323,n1324,n1325,n1326,n1327,n1328,n1329,
n1330,n1331,n1332,n1333,n1334,n1335,n1336,n1337,n1338,n1339,
n1340,n1341,n1342,n1343,n1344,n1345,n1346,n1347,n1348,n1349,
n1350,n1351,n1352,n1353,n1354,n1355,n1356,n1357,n1358,n1359,
n1360,n1361,n1362,n1363,n1364,n1365,n1366,n1367,n1368,n1369,
n1370,n1371,n1372,n1373,n1374,n1375,n1376,n1377,n1378,n1379,
n1380,n1381,n1382,n1383,n1384,n1385,n1386,n1387,n1389,n1390,
n1391,n1392,n1393,n1394,n1395,n1396,n1397,n1398,n1399,n1400,
n1401,n1402,n1403,n1404,n1405,n1406,n1407,n1408,n1409,n1410,
n1411,n1412,n1413,n1414,n1415,n1416,n1417,n1418,n1419,n1420,
n1421,n1422,n1423,n1424,n1425,n1426,n1427,n1428,n1429,n1430,
n1431,n1432,n1433,n1434,n1435,n1436,n1437,n1438,n1439,n1440,
n1441,n1442,n1443,n1444,n1445,n1446,n1447,n1448,n1449,n1450,
n1451,n1452,n1453,n1454,n1455,n1456,n1457,n1458,n1459,n1460,
n1461,n1462,n1463,n1464,n1465,n1466,n1467,n1468,n1469,n1470,
n1471,n1472,n1473,n1474,n1475,n1476,n1477,n1478,n1479,n1480,
n1481,n1482,n1483,n1484,n1485,n1486,n1487,n1488,n1489,n1490,
n1491,n1492,n1493,n1494,n1495,n1496,n1497,n1498,n1499,n1500,
n1501,n1502,n1503,n1504,n1505,n1506,n1507,n1508,n1509,n1510,
n1511,n1512,n1513,n1514,n1515,n1516,n1517,n1518,n1519,n1520,
n1521,n1522,n1523,n1524,n1525,n1526,n1527,n1528,n1529,n1530,
n1531,n1532,n1533,n1534,n1535,n1536,n1537,n1538,n1539,n1540,
n1541,n1542,n1543,n1544,n1545,n1546,n1547,n1548,n1549,n1550,
n1551,n1552,n1553,n1554,n1555,n1556,n1557,n1558,n1559,n1560,
n1561,n1562,n1563,n1564,n1565,n1566,n1567,n1568,n1569,n1570,
n1571,n1572,n1573,n1574,n1575,n1576,n1577,n1578,n1579,n1580,
n1581,n1582,n1583,n1584,n1585,n1586,n1587,n1588,n1589,n1590,
n1591,n1592,n1593,n1594,n1595,n1596,n1597,n1598,n1599,n1600,
n1601,n1602,n1603,n1604,n1605,n1606,n1607,n1608,n1609,n1610,
n1611,n1612,n1613,n1614,n1615,n1616,n1617,n1618,n1619,n1620,
n1621,n1622,n1623,n1624,n1625,n1626,n1627,n1628,n1629,n1630,
n1631,n1632,n1633,n1634,n1635,n1636,n1637,n1638,n1639,n1640,
n1641,n1642,n1643,n1644,n1645,n1646,n1647,n1648,n1649,n1650,
n1651,n1652,n1653,n1654,n1655,n1656,n1657,n1658,n1659,n1660,
n1661,n1662,n1663,n1664,n1665,n1666,n1667,n1668,n1669,n1670,
n1671,n1672,n1673,n1674,n1675,n1676,n1677,n1678,n1679,n1680,
n1681,n1682,n1683,n1684,n1685,n1686,n1687,n1688,n1689,n1690,
n1691,n1692,n1693,n1694,n1695,n1696,n1697,n1698,n1699,n1700,
n1701,n1702,n1703,n1704,n1705,n1706,n1707,n1708,n1709,n1710,
n1711,n1712,n1713,n1714,n1715,n1716,n1717,n1718,n1719,n1720,
n1721,n1722,n1723,n1724,n1725,n1726,n1727,n1728,n1729,n1730,
n1731,n1732,n1733,n1734,n1735,n1736,n1737,n1738,n1739,n1740,
n1741,n1742,n1743,n1744,n1745,n1746,n1747,n1748,n1749,n1750,
n1751,n1752,n1753,n1754,n1755,n1756,n1757,n1758,n1759,n1760,
n1761,n1762,n1763,n1764,n1765,n1766,n1767,n1768,n1769,n1770,
n1771,n1772,n1773,n1774,n1775,n1776,n1777,n1778,n1779,n1780,
n1781,n1782,n1783,n1784,n1785,n1786,n1787,n1788,n1789,n1790,
n1791,n1792,n1793,n1794,n1795,n1796,n1797,n1798,n1799,n1800,
n1801,n1802,n1803,n1804,n1805,n1806,n1807,n1808,n1809,n1810,
n1811,n1812,n1813,n1814,n1815,n1816,n1817,n1818,n1819,n1820,
n1821,n1822,n1823,n1824,n1825,n1826,n1827,n1828,n1829,n1830,
n1831,n1832,n1833,n1834,n1835,n1836,n1837,n1838,n1839,n1840,
n1841,n1842,n1843,n1844,n1845,n1846,n1847,n1848,n1849,n1850,
n1851,n1852,n1853,n1854,n1855,n1856,n1857,n1858,n1859,n1860,
n1861,n1862,n1863,n1864,n1865,n1866,n1867,n1868,n1869,n1870,
n1871,n1872,n1873,n1874,n1875,n1876,n1877,n1878,n1879,n1880,
n1881,n1882,n1883,n1884,n1885,n1886,n1887,n1888,n1889,n1890,
n1891,n1892,n1893,n1894,n1895,n1896,n1897,n1898,n1899,n1900,
n1901,n1902,n1903,n1905,n1906,n1907,n1908,n1909,n1910,n1911,
n1912,n1913,n1914,n1915,n1916,n1917,n1918,n1919,n1920,n1921,
n1922,n1923,n1924,n1925,n1926,n1927,n1928,n1929,n1930,n1931,
n1932,n1933,n1934,n1935,n1936,n1937,n1938,n1939,n1940,n1941,
n1942,n1943,n1944,n1945,n1946,n1947,n1948,n1949,n1950,n1951,
n1952,n1953,n1954,n1955,n1956,n1957,n1958,n1959,n1960,n1961,
n1962,n1963,n1964,n1965,n1966,n1967,n1968,n1969,n1970,n1971,
n1972,n1973,n1974,n1975,n1976,n1977,n1978,n1979,n1980,n1981,
n1982,n1983,n1984,n1985,n1986,n1987,n1988,n1989,n1990,n1991,
n1992,n1993,n1994,n1995,n1996,n1997,n1998,n1999,n2000,n2001,
n2002,n2003,n2004,n2005,n2006,n2007,n2008,n2009,n2010,n2011,
n2012,n2013,n2014,n2015,n2016,n2017,n2018,n2019,n2020,n2021,
n2022,n2023,n2024,n2025,n2026,n2027,n2028,n2029,n2030,n2031,
n2032,n2033,n2034,n2035,n2036,n2037,n2038,n2039,n2040,n2041,
n2042,n2043,n2044,n2045,n2046,n2047,n2048,n2049,n2050,n2051,
n2052,n2053,n2054,n2055,n2056,n2057,n2058,n2059,n2060,n2061,
n2062,n2063,n2064,n2065,n2066,n2067,n2068,n2069,n2070,n2071,
n2072,n2073,n2074,n2075,n2076,n2077,n2078,n2079,n2080,n2081,
n2082,n2083,n2084,n2085,n2086,n2087,n2088,n2089,n2090,n2091,
n2092,n2093,n2094,n2095,n2096,n2097,n2098,n2099,n2100,n2101,
n2102,n2103,n2104,n2105,n2106,n2107,n2108,n2109,n2110,n2111,
n2112,n2113,n2114,n2115,n2116,n2117,n2118,n2119,n2120,n2121,
n2122,n2123,n2124,n2125,n2126,n2127,n2128,n2129,n2130,n2131,
n2132,n2133,n2134,n2135,n2136,n2137,n2138,n2139,n2140,n2141,
n2142,n2143,n2144,n2145,n2146,n2147,n2148,n2149,n2150,n2151,
n2152,n2153,n2154,n2155,n2156,n2157,n2158,n2159,n2160,n2161,
n2162,n2163,n2164,n2165,n2166,n2167,n2168,n2169,n2170,n2171,
n2172,n2173,n2174,n2175,n2176,n2177,n2178,n2179,n2180,n2181,
n2182,n2183,n2184,n2185,n2186,n2187,n2188,n2189,n2190,n2191,
n2192,n2193,n2194,n2195,n2196,n2197,n2198,n2199,n2200,n2201,
n2202,n2203,n2204,n2205,n2206,n2207,n2208,n2209,n2210,n2211,
n2212,n2213,n2214,n2215,n2216,n2217,n2218,n2219,n2220,n2221,
n2222,n2223,n2224,n2225,n2226,n2227,n2228,n2229,n2230,n2231,
n2232,n2233,n2234,n2235,n2236,n2237,n2238,n2239,n2240,n2241,
n2242,n2243,n2244,n2245,n2246,n2247,n2248,n2249,n2250,n2251,
n2252,n2253,n2254,n2255,n2256,n2257,n2258,n2259,n2260,n2261,
n2262,n2263,n2264,n2265,n2266,n2267,n2268,n2269,n2270,n2271,
n2272,n2273,n2274,n2275,n2276,n2277,n2278,n2279,n2280,n2281,
n2282,n2283,n2284,n2285,n2286,n2287,n2288,n2289,n2290,n2291,
n2292,n2293,n2294,n2295,n2296,n2297,n2298,n2299,n2300,n2301,
n2302,n2303,n2304,n2305,n2306,n2307,n2308,n2309,n2310,n2311,
n2312,n2313,n2314,n2315,n2316,n2317,n2318,n2319,n2320,n2321,
n2322,n2323,n2324,n2325,n2326,n2327,n2328,n2329,n2330,n2331,
n2332,n2333,n2334,n2335,n2336,n2337,n2338,n2339,n2340,n2341,
n2342,n2343,n2344,n2345,n2346,n2347,n2348,n2349,n2350,n2351,
n2352,n2353,n2354,n2355,n2356,n2357,n2358,n2359,n2360,n2361,
n2362,n2363,n2364,n2365,n2366,n2367,n2368,n2369,n2370,n2371,
n2372,n2373,n2374,n2375,n2376,n2377,n2378,n2379,n2380,n2381,
n2382,n2383,n2384,n2385,n2386,n2387,n2388,n2389,n2390,n2391,
n2392,n2393,n2394,n2395,n2396,n2397,n2398,n2399,n2400,n2401,
n2402,n2403,n2404,n2405,n2406,n2407,n2408,n2409,n2410,n2411,
n2412,n2413,n2414,n2415,n2416,n2417,n2418,n2419,n2420,n2421,
n2422,n2423,n2424,n2425,n2426,n2427,n2428,n2430,n2431,n2432,
n2433,n2434,n2435,n2436,n2437,n2438,n2439,n2440,n2441,n2442,
n2443,n2444,n2445,n2446,n2447,n2448,n2449,n2450,n2451,n2452,
n2453,n2454,n2455,n2456,n2457,n2458,n2459,n2460,n2461,n2462,
n2463,n2464,n2465,n2466,n2467,n2468,n2469,n2470,n2471,n2472,
n2473,n2474,n2475,n2476,n2477,n2478,n2479,n2480,n2481,n2482,
n2483,n2484,n2485,n2486,n2487,n2488,n2489,n2490,n2491,n2492,
n2493,n2494,n2495,n2496,n2497,n2498,n2499,n2500,n2501,n2502,
n2503,n2504,n2505,n2506,n2507,n2508,n2509,n2510,n2511,n2512,
n2513,n2514,n2515,n2516,n2517,n2518,n2519,n2520,n2521,n2522,
n2523,n2524,n2525,n2526,n2527,n2528,n2529,n2530,n2531,n2532,
n2533,n2534,n2535,n2536,n2537,n2538,n2539,n2540,n2541,n2542,
n2543,n2544,n2545,n2546,n2547,n2548,n2549,n2550,n2551,n2552,
n2553,n2554,n2555,n2556,n2557,n2558,n2559,n2560,n2561,n2562,
n2563,n2564,n2565,n2566,n2567,n2568,n2569,n2570,n2571,n2572,
n2573,n2574,n2575,n2576,n2577,n2578,n2579,n2580,n2581,n2582,
n2583,n2584,n2585,n2586,n2587,n2588,n2589,n2590,n2591,n2592,
n2593,n2594,n2595,n2596,n2597,n2598,n2599,n2600,n2601,n2602,
n2603,n2604,n2605,n2606,n2607,n2608,n2609,n2610,n2611,n2612,
n2613,n2614,n2615,n2616,n2617,n2618,n2619,n2620,n2621,n2622,
n2623,n2624,n2625,n2626,n2627,n2628,n2629,n2630,n2631,n2632,
n2633,n2634,n2635,n2636,n2637,n2638,n2639,n2640,n2641,n2642,
n2643,n2644,n2645,n2646,n2647,n2648,n2649,n2650,n2651,n2652,
n2653,n2654,n2655,n2656,n2657,n2658,n2659,n2660,n2661,n2662,
n2663,n2664,n2665,n2666,n2667,n2668,n2669,n2670,n2671,n2672,
n2673,n2674,n2675,n2676,n2677,n2678,n2679,n2680,n2681,n2682,
n2683,n2684,n2685,n2686,n2687,n2688,n2689,n2690,n2691,n2692,
n2693,n2694,n2695,n2696,n2697,n2698,n2699,n2700,n2701,n2702,
n2703,n2704,n2705,n2706,n2707,n2708,n2709,n2710,n2711,n2712,
n2713,n2714,n2715,n2716,n2717,n2718,n2719,n2720,n2721,n2722,
n2723,n2724,n2725,n2726,n2727,n2728,n2729,n2730,n2731,n2732,
n2733,n2734,n2735,n2736,n2737,n2738,n2739,n2740,n2741,n2742,
n2743,n2744,n2745,n2746,n2747,n2748,n2749,n2750,n2751,n2752,
n2753,n2754,n2755,n2756,n2757,n2758,n2759,n2760,n2761,n2762,
n2763,n2764,n2765,n2766,n2767,n2768,n2769,n2770,n2771,n2772,
n2773,n2774,n2775,n2776,n2777,n2778,n2779,n2780,n2781,n2782,
n2783,n2784,n2785,n2786,n2787,n2788,n2789,n2790,n2791,n2792,
n2793,n2794,n2795,n2796,n2797,n2798,n2799,n2800,n2801,n2802,
n2803,n2804,n2805,n2806,n2807,n2808,n2809,n2810,n2811,n2812,
n2813,n2814,n2815,n2816,n2817,n2818,n2819,n2820,n2821,n2822,
n2823,n2824,n2825,n2826,n2827,n2828,n2829,n2830,n2831,n2832,
n2833,n2834,n2835,n2836,n2837,n2838,n2839,n2840,n2841,n2842,
n2843,n2844,n2845,n2846,n2847,n2848,n2849,n2850,n2851,n2852,
n2853,n2854,n2855,n2856,n2857,n2858,n2859,n2860,n2861,n2862,
n2863,n2864,n2865,n2866,n2867,n2868,n2869,n2870,n2871,n2872,
n2873,n2874,n2875,n2876,n2877,n2878,n2879,n2880,n2881,n2882,
n2883,n2884,n2885,n2886,n2887,n2888,n2889,n2890,n2891,n2893,
n2894,n2895,n2896,n2897,n2898,n2899,n2900,n2901,n2902,n2903,
n2904,n2905,n2906,n2907,n2908,n2909,n2910,n2911,n2912,n2913,
n2914,n2915,n2916,n2917,n2918,n2919,n2920,n2921,n2922,n2923,
n2924,n2925,n2926,n2927,n2928,n2929,n2930,n2931,n2932,n2933,
n2934,n2935,n2936,n2937,n2938,n2939,n2940,n2941,n2942,n2943,
n2944,n2945,n2946,n2947,n2948,n2949,n2950,n2951,n2952,n2953,
n2954,n2955,n2956,n2957,n2958,n2959,n2960,n2961,n2962,n2963,
n2964,n2965,n2966,n2967,n2968,n2969,n2970,n2971,n2972,n2973,
n2974,n2975,n2976,n2977,n2978,n2979,n2980,n2981,n2982,n2983,
n2984,n2985,n2986,n2987,n2988,n2989,n2990,n2991,n2992,n2993,
n2994,n2995,n2996,n2997,n2998,n2999,n3000,n3001,n3002,n3003,
n3004,n3005,n3006,n3007,n3008,n3009,n3010,n3011,n3012,n3013,
n3014,n3015,n3016,n3017,n3018,n3019,n3020,n3021,n3022,n3023,
n3024,n3025,n3026,n3027,n3028,n3029,n3030,n3031,n3032,n3033,
n3034,n3035,n3036,n3037,n3038,n3039,n3040,n3041,n3042,n3043,
n3044,n3045,n3046,n3047,n3048,n3049,n3050,n3051,n3052,n3053,
n3054,n3055,n3056,n3057,n3058,n3059,n3060,n3061,n3062,n3063,
n3064,n3065,n3066,n3067,n3068,n3069,n3070,n3071,n3072,n3073,
n3074,n3075,n3076,n3077,n3078,n3079,n3080,n3081,n3082,n3083,
n3084,n3085,n3086,n3087,n3088,n3089,n3090,n3091,n3092,n3093,
n3094,n3095,n3096,n3097,n3098,n3099,n3100,n3101,n3102,n3103,
n3104,n3105,n3106,n3107,n3108,n3109,n3110,n3111,n3112,n3113,
n3114,n3115,n3116,n3117,n3118,n3119,n3120,n3121,n3122,n3123,
n3124,n3125,n3126,n3127,n3128,n3129,n3130,n3131,n3132,n3133,
n3134,n3135,n3136,n3137,n3138,n3139,n3140,n3141,n3142,n3143,
n3144,n3145,n3146,n3147,n3148,n3149,n3150,n3151,n3152,n3153,
n3154,n3155,n3156,n3157,n3158,n3159,n3160,n3161,n3162,n3163,
n3164,n3165,n3166,n3167,n3168,n3169,n3170,n3171,n3172,n3173,
n3174,n3175,n3176,n3177,n3178,n3179,n3180,n3181,n3182,n3183,
n3184,n3185,n3186,n3187,n3188,n3189,n3190,n3191,n3192,n3193,
n3194,n3195,n3196,n3197,n3198,n3199,n3200,n3201,n3202,n3203,
n3204,n3205,n3206,n3207,n3208,n3209,n3210,n3211,n3212,n3213,
n3214,n3215,n3216,n3217,n3218,n3219,n3220,n3221,n3222,n3223,
n3224,n3225,n3226,n3227,n3228,n3229,n3230,n3231,n3232,n3233,
n3234,n3235,n3236,n3237,n3238,n3239,n3240,n3241,n3242,n3243,
n3244,n3245,n3246,n3247,n3248,n3249,n3250,n3251,n3252,n3253,
n3254,n3255,n3256,n3257,n3258,n3259,n3260,n3261,n3262,n3263,
n3264,n3265,n3266,n3267,n3268,n3269,n3270,n3271,n3272,n3273,
n3274,n3275,n3276,n3277,n3278,n3279,n3280,n3281,n3282,n3283,
n3284,n3285,n3286,n3287,n3288,n3289,n3290,n3291,n3292,n3293,
n3294,n3295,n3296,n3297,n3298,n3299,n3300,n3301,n3302,n3303,
n3304,n3305,n3306,n3307,n3308,n3309,n3310,n3311,n3312,n3313,
n3314,n3315,n3316,n3317,n3318,n3319,n3320,n3321,n3322,n3323,
n3324,n3325,n3326,n3327,n3328,n3329,n3330,n3331,n3332,n3333,
n3334,n3335,n3336,n3337,n3338,n3339,n3340,n3341,n3342,n3343,
n3344,n3345,n3346,n3347,n3348,n3349,n3350,n3351,n3352,n3354,
n3355,n3356,n3357,n3358,n3359,n3360,n3361,n3362,n3363,n3364,
n3365,n3366,n3367,n3368,n3369,n3370,n3371,n3372,n3373,n3374,
n3375,n3376,n3377,n3378,n3379,n3380,n3381,n3382,n3383,n3384,
n3385,n3386,n3387,n3388,n3389,n3390,n3391,n3392,n3393,n3394,
n3395,n3396,n3397,n3398,n3399,n3400,n3401,n3402,n3403,n3404,
n3405,n3406,n3407,n3408,n3409,n3410,n3411,n3412,n3413,n3414,
n3415,n3416,n3417,n3418,n3419,n3420,n3421,n3422,n3423,n3424,
n3425,n3426,n3427,n3428,n3429,n3430,n3431,n3432,n3433,n3434,
n3435,n3436,n3437,n3438,n3439,n3440,n3441,n3442,n3443,n3444,
n3445,n3446,n3447,n3448,n3449,n3450,n3451,n3452,n3453,n3454,
n3455,n3456,n3457,n3458,n3459,n3460,n3461,n3462,n3463,n3464,
n3465,n3466,n3467,n3468,n3469,n3470,n3471,n3472,n3473,n3474,
n3475,n3476,n3477,n3478,n3479,n3480,n3481,n3482,n3483,n3484,
n3485,n3486,n3487,n3488,n3489,n3490,n3491,n3492,n3493,n3494,
n3495,n3496,n3497,n3498,n3499,n3500,n3501,n3502,n3503,n3504,
n3505,n3506,n3507,n3508,n3509,n3510,n3511,n3512,n3513,n3514,
n3515,n3516,n3517,n3518,n3519,n3520,n3521,n3522,n3523,n3524,
n3525,n3526,n3527,n3528,n3529,n3530,n3531,n3532,n3533,n3534,
n3535,n3536,n3537,n3538,n3539,n3540,n3541,n3542,n3543,n3544,
n3545,n3546,n3547,n3548,n3549,n3550,n3551,n3552,n3553,n3554,
n3555,n3556,n3557,n3558,n3559,n3560,n3561,n3562,n3563,n3564,
n3565,n3566,n3567,n3568,n3569,n3570,n3571,n3572,n3573,n3574,
n3575,n3576,n3577,n3578,n3579,n3580,n3581,n3582,n3583,n3584,
n3585,n3586,n3587,n3588,n3589,n3590,n3591,n3592,n3593,n3594,
n3595,n3596,n3597,n3598,n3599,n3600,n3601,n3602,n3603,n3604,
n3605,n3606,n3607,n3608,n3609,n3610,n3611,n3612,n3613,n3614,
n3615,n3616,n3617,n3618,n3619,n3620,n3621,n3622,n3623,n3624,
n3625,n3626,n3627,n3628,n3629,n3630,n3631,n3632,n3633,n3634,
n3635,n3636,n3637,n3638,n3639,n3640,n3641,n3642,n3643,n3644,
n3645,n3646,n3647,n3648,n3649,n3650,n3651,n3652,n3653,n3654,
n3655,n3656,n3657,n3658,n3659,n3660,n3661,n3662,n3663,n3664,
n3665,n3666,n3667,n3668,n3669,n3670,n3671,n3672,n3673,n3674,
n3675,n3676,n3677,n3678,n3679,n3680,n3681,n3682,n3683,n3684,
n3685,n3686,n3687,n3688,n3689,n3690,n3691,n3692,n3693,n3694,
n3695,n3696,n3697,n3698,n3699,n3700,n3701,n3702,n3703,n3704,
n3705,n3706,n3707,n3708,n3709,n3710,n3711,n3712,n3713,n3714,
n3715,n3716,n3717,n3718,n3719,n3720,n3721,n3722,n3723,n3724,
n3725,n3726,n3727,n3728,n3729,n3730,n3731,n3732,n3733,n3734,
n3735,n3736,n3737,n3738,n3739,n3740,n3741,n3742,n3743,n3744,
n3745,n3746,n3747,n3748,n3749,n3750,n3751,n3752,n3753,n3754,
n3755,n3756,n3757,n3758,n3759,n3760,n3761,n3762,n3763,n3764,
n3765,n3766,n3767,n3768,n3769,n3770,n3771,n3772,n3773,n3774,
n3775,n3776,n3777,n3778,n3779,n3780,n3781,n3782,n3783,n3784,
n3785,n3786,n3787,n3788,n3789,n3790,n3791,n3792,n3793,n3794,
n3795,n3796,n3797,n3798,n3799,n3800,n3801,n3802,n3803,n3804,
n3805,n3806,n3807,n3808,n3809,n3810,n3811,n3812,n3814,n3815,
n3816,n3817,n3818,n3819,n3820,n3821,n3822,n3823,n3824,n3825,
n3826,n3827,n3828,n3829,n3830,n3831,n3832,n3833,n3834,n3835,
n3836,n3837,n3838,n3839,n3840,n3841,n3842,n3843,n3844,n3845,
n3846,n3847,n3848,n3849,n3850,n3851,n3852,n3853,n3854,n3855,
n3856,n3857,n3858,n3859,n3860,n3861,n3862,n3863,n3864,n3865,
n3866,n3867,n3868,n3869,n3870,n3871,n3872,n3873,n3874,n3875,
n3876,n3877,n3878,n3879,n3880,n3881,n3882,n3883,n3884,n3885,
n3886,n3887,n3888,n3889,n3890,n3891,n3892,n3893,n3894,n3895,
n3896,n3897,n3898,n3899,n3900,n3901,n3902,n3903,n3904,n3905,
n3906,n3907,n3908,n3909,n3910,n3911,n3912,n3913,n3914,n3915,
n3916,n3917,n3918,n3919,n3920,n3921,n3922,n3923,n3924,n3925,
n3926,n3927,n3928,n3929,n3930,n3931,n3932,n3933,n3934,n3935,
n3936,n3937,n3938,n3939,n3940,n3941,n3942,n3943,n3944,n3945,
n3946,n3947,n3948,n3949,n3950,n3951,n3952,n3953,n3954,n3955,
n3956,n3957,n3958,n3959,n3960,n3961,n3962,n3963,n3964,n3965,
n3966,n3967,n3968,n3969,n3970,n3971,n3972,n3973,n3974,n3975,
n3976,n3977,n3978,n3979,n3980,n3981,n3982,n3983,n3984,n3985,
n3986,n3987,n3988,n3989,n3990,n3991,n3992,n3993,n3994,n3995,
n3996,n3997,n3998,n3999,n4000,n4001,n4002,n4003,n4004,n4005,
n4006,n4007,n4008,n4009,n4010,n4011,n4012,n4013,n4014,n4015,
n4016,n4017,n4018,n4019,n4020,n4021,n4022,n4023,n4024,n4025,
n4026,n4027,n4028,n4029,n4030,n4031,n4032,n4033,n4034,n4035,
n4036,n4037,n4038,n4039,n4040,n4041,n4042,n4043,n4044,n4045,
n4046,n4047,n4048,n4049,n4050,n4051,n4052,n4053,n4054,n4055,
n4056,n4057,n4058,n4059,n4060,n4061,n4062,n4063,n4064,n4065,
n4066,n4067,n4068,n4069,n4070,n4071,n4072,n4073,n4074,n4075,
n4076,n4077,n4078,n4079,n4080,n4081,n4082,n4083,n4084,n4085,
n4086,n4087,n4088,n4089,n4090,n4091,n4092,n4093,n4094,n4095,
n4096,n4097,n4098,n4099,n4100,n4101,n4102,n4103,n4104,n4105,
n4106,n4107,n4108,n4109,n4110,n4111,n4112,n4113,n4114,n4115,
n4116,n4117,n4118,n4119,n4120,n4121,n4122,n4123,n4124,n4125,
n4126,n4127,n4128,n4129,n4130,n4131,n4132,n4133,n4134,n4135,
n4136,n4137,n4138,n4139,n4140,n4141,n4142,n4143,n4144,n4145,
n4146,n4147,n4148,n4149,n4150,n4151,n4152,n4153,n4154,n4155,
n4156,n4157,n4158,n4159,n4160,n4161,n4162,n4163,n4164,n4165,
n4166,n4167,n4168,n4169,n4170,n4171,n4172,n4173,n4174,n4175,
n4176,n4177,n4178,n4179,n4180,n4181,n4182,n4183,n4184,n4185,
n4186,n4187,n4188,n4189,n4190,n4191,n4192,n4193,n4194,n4195,
n4196,n4197,n4198,n4199,n4200,n4201,n4202,n4203,n4204,n4205,
n4206,n4207,n4208,n4209,n4210,n4211,n4212,n4214,n4215,n4216,
n4217,n4218,n4219,n4220,n4221,n4222,n4223,n4224,n4225,n4226,
n4227,n4228,n4229,n4230,n4231,n4232,n4233,n4234,n4235,n4236,
n4237,n4238,n4239,n4240,n4241,n4242,n4243,n4244,n4245,n4246,
n4247,n4248,n4249,n4250,n4251,n4252,n4253,n4254,n4255,n4256,
n4257,n4258,n4259,n4260,n4261,n4262,n4263,n4264,n4265,n4266,
n4267,n4268,n4269,n4270,n4271,n4272,n4273,n4274,n4275,n4276,
n4277,n4278,n4279,n4280,n4281,n4282,n4283,n4284,n4285,n4286,
n4287,n4288,n4289,n4290,n4291,n4292,n4293,n4294,n4295,n4296,
n4297,n4298,n4299,n4300,n4301,n4302,n4303,n4304,n4305,n4306,
n4307,n4308,n4309,n4310,n4311,n4312,n4313,n4314,n4315,n4316,
n4317,n4318,n4319,n4320,n4321,n4322,n4323,n4324,n4325,n4326,
n4327,n4328,n4329,n4330,n4331,n4332,n4333,n4334,n4335,n4336,
n4337,n4338,n4339,n4340,n4341,n4342,n4343,n4344,n4345,n4346,
n4347,n4348,n4349,n4350,n4351,n4352,n4353,n4354,n4355,n4356,
n4357,n4358,n4359,n4360,n4361,n4362,n4363,n4364,n4365,n4366,
n4367,n4368,n4369,n4370,n4371,n4372,n4373,n4374,n4375,n4376,
n4377,n4378,n4379,n4380,n4381,n4382,n4383,n4384,n4385,n4386,
n4387,n4388,n4389,n4390,n4391,n4392,n4393,n4394,n4395,n4396,
n4397,n4398,n4399,n4400,n4401,n4402,n4403,n4404,n4405,n4406,
n4407,n4408,n4409,n4410,n4411,n4412,n4413,n4414,n4415,n4416,
n4417,n4418,n4419,n4420,n4421,n4422,n4423,n4424,n4425,n4426,
n4427,n4428,n4429,n4430,n4431,n4432,n4433,n4434,n4435,n4436,
n4437,n4438,n4439,n4440,n4441,n4442,n4443,n4444,n4445,n4446,
n4447,n4448,n4449,n4450,n4451,n4452,n4453,n4454,n4455,n4456,
n4457,n4458,n4459,n4460,n4461,n4462,n4463,n4464,n4465,n4466,
n4467,n4468,n4469,n4470,n4471,n4472,n4473,n4474,n4475,n4476,
n4477,n4478,n4479,n4480,n4481,n4482,n4483,n4484,n4485,n4486,
n4487,n4488,n4489,n4490,n4491,n4492,n4493,n4494,n4495,n4496,
n4497,n4498,n4499,n4500,n4501,n4502,n4503,n4504,n4505,n4506,
n4507,n4508,n4509,n4510,n4511,n4512,n4513,n4514,n4515,n4516,
n4517,n4518,n4519,n4520,n4521,n4522,n4523,n4524,n4525,n4526,
n4527,n4528,n4529,n4530,n4531,n4532,n4533,n4534,n4535,n4536,
n4537,n4538,n4539,n4540,n4541,n4542,n4543,n4544,n4545,n4546,
n4547,n4548,n4549,n4550,n4551,n4552,n4553,n4554,n4555,n4556,
n4557,n4558,n4559,n4560,n4561,n4562,n4563,n4564,n4565,n4566,
n4567,n4568,n4569,n4570,n4571,n4572,n4573,n4574,n4575,n4576,
n4577,n4578,n4579,n4580,n4581,n4582,n4583,n4584,n4585,n4586,
n4587,n4588,n4589,n4590,n4591,n4592,n4593,n4594,n4595,n4596,
n4597,n4598,n4599,n4600,n4601,n4602,n4603,n4604,n4605,n4606,
n4607,n4608,n4609,n4610,n4611,n4612,n4613,n4614,n4615,n4616,
n4617,n4618,n4619,n4620,n4621,n4622,n4623,n4624,n4625,n4626,
n4627,n4628,n4629,n4630,n4631,n4632,n4633,n4634,n4635,n4636,
n4637,n4638,n4639,n4640,n4641,n4642,n4643,n4644,n4645,n4646,
n4647,n4648,n4649,n4650,n4651,n4652,n4653,n4654,n4655,n4656,
n4657,n4659,n4660,n4661,n4662,n4663,n4664,n4665,n4666,n4667,
n4668,n4669,n4670,n4671,n4672,n4673,n4674,n4675,n4676,n4677,
n4678,n4679,n4680,n4681,n4682,n4683,n4684,n4685,n4686,n4687,
n4688,n4689,n4690,n4691,n4692,n4693,n4694,n4695,n4696,n4697,
n4698,n4699,n4700,n4701,n4702,n4703,n4704,n4705,n4706,n4707,
n4708,n4709,n4710,n4711,n4712,n4713,n4714,n4715,n4716,n4717,
n4718,n4719,n4720,n4721,n4722,n4723,n4724,n4725,n4726,n4727,
n4728,n4729,n4730,n4731,n4732,n4733,n4734,n4735,n4736,n4737,
n4738,n4739,n4740,n4741,n4742,n4743,n4744,n4745,n4746,n4747,
n4748,n4749,n4750,n4751,n4752,n4753,n4754,n4755,n4756,n4757,
n4758,n4759,n4760,n4761,n4762,n4763,n4764,n4765,n4766,n4767,
n4768,n4769,n4770,n4771,n4772,n4773,n4774,n4775,n4776,n4777,
n4778,n4779,n4780,n4781,n4782,n4783,n4784,n4785,n4786,n4787,
n4788,n4789,n4790,n4791,n4792,n4793,n4794,n4795,n4796,n4797,
n4798,n4799,n4800,n4801,n4802,n4803,n4804,n4805,n4806,n4807,
n4808,n4809,n4810,n4811,n4812,n4813,n4814,n4815,n4816,n4817,
n4818,n4819,n4820,n4821,n4822,n4823,n4824,n4825,n4826,n4827,
n4828,n4829,n4830,n4831,n4832,n4833,n4834,n4835,n4836,n4837,
n4838,n4839,n4840,n4841,n4842,n4843,n4844,n4845,n4846,n4847,
n4848,n4849,n4850,n4851,n4852,n4853,n4854,n4855,n4856,n4857,
n4858,n4859,n4860,n4861,n4862,n4863,n4864,n4865,n4866,n4867,
n4868,n4869,n4870,n4871,n4872,n4873,n4874,n4875,n4876,n4877,
n4878,n4879,n4880,n4881,n4882,n4883,n4884,n4885,n4886,n4887,
n4888,n4889,n4890,n4891,n4892,n4893,n4894,n4895,n4896,n4897,
n4898,n4899,n4900,n4901,n4902,n4903,n4904,n4905,n4906,n4907,
n4908,n4909,n4910,n4911,n4912,n4913,n4914,n4915,n4916,n4917,
n4918,n4919,n4920,n4921,n4922,n4923,n4924,n4925,n4926,n4927,
n4928,n4929,n4930,n4931,n4932,n4933,n4934,n4935,n4936,n4937,
n4938,n4939,n4940,n4941,n4942,n4943,n4944,n4945,n4946,n4947,
n4948,n4949,n4950,n4951,n4952,n4953,n4954,n4955,n4956,n4957,
n4958,n4959,n4960,n4961,n4962,n4963,n4964,n4965,n4966,n4967,
n4968,n4969,n4970,n4971,n4972,n4973,n4974,n4975,n4976,n4977,
n4978,n4979,n4980,n4981,n4982,n4983,n4984,n4985,n4986,n4987,
n4988,n4989,n4990,n4991,n4992,n4993,n4994,n4995,n4996,n4997,
n4998,n4999,n5000,n5001,n5002,n5003,n5004,n5005,n5006,n5007,
n5008,n5009,n5010,n5011,n5012,n5013,n5014,n5015,n5016,n5017,
n5018,n5019,n5020,n5021,n5022,n5023,n5024,n5025,n5026,n5027,
n5028,n5029,n5030,n5031,n5032,n5033,n5034,n5035,n5036,n5037,
n5038,n5039,n5040,n5041,n5042,n5043,n5044,n5045,n5046,n5047,
n5048,n5049,n5050,n5051,n5052,n5053,n5054,n5055,n5056,n5057,
n5058,n5059,n5060,n5061,n5062,n5063,n5064,n5065,n5066,n5067,
n5068,n5069,n5070,n5071,n5072,n5073,n5074,n5075,n5076,n5077,
n5078,n5079,n5080,n5081,n5082,n5083,n5084;
not gate_0(n20,pi0);
not gate_1(n21,pi1);
not gate_2(n22,pi2);
not gate_3(n23,pi3);
not gate_4(n24,pi4);
not gate_5(n25,pi5);
not gate_6(n26,pi6);
not gate_7(n27,pi7);
not gate_8(n28,pi8);
not gate_9(n29,pi9);
and gate_10(n30,pi2,pi3);
not gate_11(n31,n30);
and gate_12(n32,n28,pi9);
not gate_13(n33,n32);
and gate_14(n34,pi6,n32);
and gate_15(n35,n30,n34);
not gate_16(n36,n35);
and gate_17(n37,n22,n23);
not gate_18(n38,n37);
and gate_19(n39,pi8,n29);
not gate_20(n40,n39);
and gate_21(n41,n26,n39);
not gate_22(n42,n41);
and gate_23(n43,n37,n41);
not gate_24(n44,n43);
and gate_25(n45,n36,n44);
not gate_26(n46,n45);
and gate_27(n47,n20,n21);
not gate_28(n48,n47);
and gate_29(n49,n25,pi7);
not gate_30(n50,n49);
and gate_31(n51,pi4,n49);
not gate_32(n52,n51);
and gate_33(n53,n47,n51);
not gate_34(n54,n53);
and gate_35(n55,pi0,pi1);
and gate_36(n56,pi5,n27);
not gate_37(n57,n56);
and gate_38(n58,n24,n56);
not gate_39(n59,n58);
and gate_40(n60,n55,n58);
not gate_41(n61,n60);
and gate_42(n62,n54,n61);
not gate_43(n63,n62);
and gate_44(n64,n46,n63);
not gate_45(n65,n64);
and gate_46(n66,pi1,pi2);
not gate_47(n67,n66);
and gate_48(n68,n20,n66);
and gate_49(n69,n25,n26);
not gate_50(n70,n69);
and gate_51(n71,n24,n69);
and gate_52(n72,n68,n71);
not gate_53(n73,n72);
and gate_54(n74,n22,pi4);
not gate_55(n75,n74);
and gate_56(n76,n20,pi1);
not gate_57(n77,n76);
and gate_58(n78,n74,n76);
not gate_59(n79,n78);
and gate_60(n80,pi2,n24);
not gate_61(n81,n80);
and gate_62(n82,n75,n81);
not gate_63(n83,n82);
and gate_64(n84,pi0,n21);
not gate_65(n85,n84);
and gate_66(n86,n83,n84);
not gate_67(n87,n86);
and gate_68(n88,n79,n87);
not gate_69(n89,n88);
and gate_70(n90,pi5,pi6);
not gate_71(n91,n90);
and gate_72(n92,n89,n90);
not gate_73(n93,n92);
and gate_74(n94,n73,n93);
not gate_75(n95,n94);
and gate_76(n96,pi9,n95);
not gate_77(n97,n96);
and gate_78(n98,pi1,n24);
and gate_79(n99,n25,pi6);
not gate_80(n100,n99);
and gate_81(n101,n22,n99);
and gate_82(n102,n98,n101);
not gate_83(n103,n102);
and gate_84(n104,n21,pi2);
not gate_85(n105,n104);
and gate_86(n106,pi4,n26);
not gate_87(n107,n106);
and gate_88(n108,n104,n106);
not gate_89(n109,n108);
and gate_90(n110,pi5,n108);
not gate_91(n111,n110);
and gate_92(n112,n103,n111);
not gate_93(n113,n112);
and gate_94(n114,pi0,n29);
and gate_95(n115,n113,n114);
not gate_96(n116,n115);
and gate_97(n117,n97,n116);
not gate_98(n118,n117);
and gate_99(n119,n27,n118);
not gate_100(n120,n119);
and gate_101(n121,pi5,n29);
not gate_102(n122,n121);
and gate_103(n123,pi6,pi9);
not gate_104(n124,n123);
and gate_105(n125,n25,n123);
not gate_106(n126,n125);
and gate_107(n127,n122,n126);
not gate_108(n128,n127);
and gate_109(n129,pi2,n128);
not gate_110(n130,n129);
and gate_111(n131,n22,n25);
not gate_112(n132,n131);
and gate_113(n133,n26,n29);
not gate_114(n134,n133);
and gate_115(n135,n131,n133);
not gate_116(n136,n135);
and gate_117(n137,n130,n136);
not gate_118(n138,n137);
and gate_119(n139,pi4,pi7);
not gate_120(n140,n139);
and gate_121(n141,n21,n139);
and gate_122(n142,n138,n141);
and gate_123(n143,pi0,n142);
not gate_124(n144,n143);
and gate_125(n145,n120,n144);
not gate_126(n146,n145);
and gate_127(n147,n23,n146);
not gate_128(n148,n147);
and gate_129(n149,pi5,pi7);
not gate_130(n150,n149);
and gate_131(n151,n80,n149);
not gate_132(n152,n151);
and gate_133(n153,n25,n27);
not gate_134(n154,n153);
and gate_135(n155,n74,n153);
not gate_136(n156,n155);
and gate_137(n157,n152,n156);
not gate_138(n158,n157);
and gate_139(n159,n20,n26);
not gate_140(n160,n159);
and gate_141(n161,n158,n159);
not gate_142(n162,n161);
and gate_143(n163,pi0,pi5);
not gate_144(n164,n163);
and gate_145(n165,n22,n24);
and gate_146(n166,pi6,n27);
not gate_147(n167,n166);
and gate_148(n168,n165,n166);
and gate_149(n169,n163,n168);
not gate_150(n170,n169);
and gate_151(n171,n162,n170);
not gate_152(n172,n171);
and gate_153(n173,pi3,n29);
not gate_154(n174,n173);
and gate_155(n175,n172,n173);
and gate_156(n176,n21,n175);
not gate_157(n177,n176);
and gate_158(n178,n148,n177);
and gate_159(n179,pi7,pi9);
not gate_160(n180,n179);
and gate_161(n181,n27,n29);
not gate_162(n182,n181);
and gate_163(n183,n180,n182);
not gate_164(n184,n183);
and gate_165(n185,pi8,n184);
and gate_166(n186,n25,n185);
not gate_167(n187,n186);
and gate_168(n188,n27,pi9);
not gate_169(n189,n188);
and gate_170(n190,pi7,n29);
not gate_171(n191,n190);
and gate_172(n192,n189,n191);
not gate_173(n193,n192);
and gate_174(n194,n33,n40);
not gate_175(n195,n194);
and gate_176(n196,pi5,n195);
and gate_177(n197,n192,n196);
not gate_178(n198,n197);
and gate_179(n199,n187,n198);
not gate_180(n200,n199);
and gate_181(n201,n21,n200);
not gate_182(n202,n201);
and gate_183(n203,n25,n28);
not gate_184(n204,n203);
and gate_185(n205,pi5,pi8);
not gate_186(n206,n205);
and gate_187(n207,n204,n206);
not gate_188(n208,n207);
and gate_189(n209,pi7,n207);
not gate_190(n210,n209);
and gate_191(n211,pi5,n28);
not gate_192(n212,n211);
and gate_193(n213,n180,n212);
not gate_194(n214,n213);
and gate_195(n215,n210,n214);
and gate_196(n216,pi1,n215);
not gate_197(n217,n216);
and gate_198(n218,n202,n217);
not gate_199(n219,n218);
and gate_200(n220,pi3,n219);
not gate_201(n221,n220);
and gate_202(n222,n150,n154);
not gate_203(n223,n222);
and gate_204(n224,pi1,n223);
not gate_205(n225,n224);
and gate_206(n226,n21,n49);
not gate_207(n227,n226);
and gate_208(n228,n225,n227);
not gate_209(n229,n228);
and gate_210(n230,pi8,n229);
not gate_211(n231,n230);
and gate_212(n232,n27,n28);
not gate_213(n233,n232);
and gate_214(n234,n21,pi5);
and gate_215(n235,n232,n234);
not gate_216(n236,n235);
and gate_217(n237,n231,n236);
not gate_218(n238,n237);
and gate_219(n239,n23,pi9);
not gate_220(n240,n239);
and gate_221(n241,n238,n239);
not gate_222(n242,n241);
and gate_223(n243,n221,n242);
not gate_224(n244,n243);
and gate_225(n245,pi2,n244);
not gate_226(n246,n245);
and gate_227(n247,n28,n29);
not gate_228(n248,n247);
and gate_229(n249,n153,n247);
not gate_230(n250,n249);
and gate_231(n251,n198,n250);
not gate_232(n252,n251);
and gate_233(n253,pi3,n252);
not gate_234(n254,n253);
and gate_235(n255,n23,pi7);
not gate_236(n256,n255);
and gate_237(n257,n194,n212);
and gate_238(n258,n255,n257);
not gate_239(n259,n258);
and gate_240(n260,n254,n259);
not gate_241(n261,n260);
and gate_242(n262,pi1,n261);
not gate_243(n263,n262);
and gate_244(n264,pi3,n25);
not gate_245(n265,n264);
and gate_246(n266,n21,n264);
and gate_247(n267,n27,n247);
and gate_248(n268,n266,n267);
not gate_249(n269,n268);
and gate_250(n270,n263,n269);
not gate_251(n271,n270);
and gate_252(n272,n22,n271);
not gate_253(n273,n272);
and gate_254(n274,n246,n273);
not gate_255(n275,n274);
and gate_256(n276,pi4,n275);
not gate_257(n277,n276);
and gate_258(n278,pi8,pi9);
not gate_259(n279,n278);
and gate_260(n280,n23,n278);
not gate_261(n281,n280);
and gate_262(n282,pi3,n247);
not gate_263(n283,n282);
and gate_264(n284,n281,n283);
not gate_265(n285,n284);
and gate_266(n286,pi2,n285);
not gate_267(n287,n286);
and gate_268(n288,n22,pi3);
not gate_269(n289,n288);
and gate_270(n290,n278,n288);
not gate_271(n291,n290);
and gate_272(n292,n287,n291);
not gate_273(n293,n292);
and gate_274(n294,n21,n293);
not gate_275(n295,n294);
and gate_276(n296,n23,n39);
not gate_277(n297,n296);
and gate_278(n298,n66,n296);
not gate_279(n299,n298);
and gate_280(n300,n295,n299);
not gate_281(n301,n300);
and gate_282(n302,n223,n301);
not gate_283(n303,n302);
and gate_284(n304,n23,pi5);
not gate_285(n305,n304);
and gate_286(n306,n21,n304);
and gate_287(n307,n27,n278);
and gate_288(n308,n306,n307);
not gate_289(n309,n308);
and gate_290(n310,pi1,n264);
and gate_291(n311,pi7,n247);
not gate_292(n312,n311);
and gate_293(n313,n310,n311);
not gate_294(n314,n313);
and gate_295(n315,n309,n314);
not gate_296(n316,n315);
and gate_297(n317,pi2,n316);
not gate_298(n318,n317);
and gate_299(n319,pi5,n188);
not gate_300(n320,n319);
and gate_301(n321,n25,n190);
not gate_302(n322,n321);
and gate_303(n323,n320,n322);
not gate_304(n324,n323);
and gate_305(n325,pi3,pi8);
not gate_306(n326,n325);
and gate_307(n327,n23,n28);
not gate_308(n328,n327);
and gate_309(n329,n326,n328);
not gate_310(n330,n329);
and gate_311(n331,n324,n330);
not gate_312(n332,n331);
and gate_313(n333,n185,n304);
not gate_314(n334,n333);
and gate_315(n335,n332,n334);
not gate_316(n336,n335);
and gate_317(n337,n21,n22);
not gate_318(n338,n337);
and gate_319(n339,n336,n337);
not gate_320(n340,n339);
and gate_321(n341,n318,n340);
and gate_322(n342,n303,n341);
not gate_323(n343,n342);
and gate_324(n344,n24,n343);
not gate_325(n345,n344);
and gate_326(n346,n277,n345);
not gate_327(n347,n346);
and gate_328(n348,pi0,n347);
not gate_329(n349,n348);
and gate_330(n350,n21,n25);
not gate_331(n351,n350);
and gate_332(n352,n23,pi8);
not gate_333(n353,n352);
and gate_334(n354,pi3,n28);
not gate_335(n355,n354);
and gate_336(n356,n353,n355);
not gate_337(n357,n356);
and gate_338(n358,n22,n27);
not gate_339(n359,n358);
and gate_340(n360,pi2,pi7);
not gate_341(n361,n360);
and gate_342(n362,n359,n361);
not gate_343(n363,n362);
and gate_344(n364,n31,n38);
not gate_345(n365,n364);
and gate_346(n366,n362,n364);
and gate_347(n367,n357,n366);
and gate_348(n368,n350,n367);
not gate_349(n369,n368);
and gate_350(n370,pi1,pi5);
not gate_351(n371,n370);
and gate_352(n372,pi7,pi8);
not gate_353(n373,n372);
and gate_354(n374,n288,n372);
not gate_355(n375,n374);
and gate_356(n376,n370,n374);
not gate_357(n377,n376);
and gate_358(n378,n369,n377);
not gate_359(n379,n378);
and gate_360(n380,n24,pi9);
not gate_361(n381,n380);
and gate_362(n382,pi4,n29);
not gate_363(n383,n382);
and gate_364(n384,n381,n383);
not gate_365(n385,n384);
and gate_366(n386,n379,n385);
not gate_367(n387,n386);
and gate_368(n388,n30,n190);
not gate_369(n389,n388);
and gate_370(n390,n27,n289);
not gate_371(n391,n390);
and gate_372(n392,pi7,n288);
not gate_373(n393,n392);
and gate_374(n394,n391,n393);
and gate_375(n395,pi9,n394);
and gate_376(n396,n25,n395);
not gate_377(n397,n396);
and gate_378(n398,n389,n397);
and gate_379(n399,n37,n188);
and gate_380(n400,pi5,n399);
not gate_381(n401,n400);
and gate_382(n402,n398,n401);
not gate_383(n403,n402);
and gate_384(n404,pi8,n403);
not gate_385(n405,n404);
and gate_386(n406,n23,n193);
not gate_387(n407,n406);
and gate_388(n408,pi3,n179);
not gate_389(n409,n408);
and gate_390(n410,n407,n409);
not gate_391(n411,n410);
and gate_392(n412,n211,n411);
and gate_393(n413,pi2,n412);
not gate_394(n414,n413);
and gate_395(n415,n405,n414);
not gate_396(n416,n415);
and gate_397(n417,n21,n416);
not gate_398(n418,n417);
and gate_399(n419,pi7,n28);
not gate_400(n420,n419);
and gate_401(n421,n27,pi8);
not gate_402(n422,n421);
and gate_403(n423,n420,n422);
not gate_404(n424,n423);
and gate_405(n425,n50,n57);
not gate_406(n426,n425);
and gate_407(n427,pi3,n426);
and gate_408(n428,n423,n427);
not gate_409(n429,n428);
and gate_410(n430,n327,n426);
not gate_411(n431,n430);
and gate_412(n432,n429,n431);
not gate_413(n433,n432);
and gate_414(n434,pi9,n433);
not gate_415(n435,n434);
and gate_416(n436,n304,n311);
not gate_417(n437,n436);
and gate_418(n438,n435,n437);
not gate_419(n439,n438);
and gate_420(n440,n22,n439);
not gate_421(n441,n440);
and gate_422(n442,n25,n195);
not gate_423(n443,n442);
and gate_424(n444,pi5,n247);
not gate_425(n445,n444);
and gate_426(n446,n443,n445);
not gate_427(n447,n446);
and gate_428(n448,n23,n27);
not gate_429(n449,n448);
and gate_430(n450,n447,n448);
and gate_431(n451,pi2,n450);
not gate_432(n452,n451);
and gate_433(n453,n441,n452);
not gate_434(n454,n453);
and gate_435(n455,pi1,n454);
not gate_436(n456,n455);
and gate_437(n457,n418,n456);
not gate_438(n458,n457);
and gate_439(n459,pi4,n458);
not gate_440(n460,n459);
and gate_441(n461,n248,n279);
not gate_442(n462,n461);
and gate_443(n463,pi2,pi5);
not gate_444(n464,n463);
and gate_445(n465,n132,n464);
not gate_446(n466,n465);
and gate_447(n467,n462,n466);
and gate_448(n468,n23,n467);
not gate_449(n469,n468);
and gate_450(n470,pi3,n203);
and gate_451(n471,n22,n470);
not gate_452(n472,n471);
and gate_453(n473,n469,n472);
not gate_454(n474,n473);
and gate_455(n475,pi7,n474);
not gate_456(n476,n475);
and gate_457(n477,n25,n32);
not gate_458(n478,n477);
and gate_459(n479,n37,n477);
not gate_460(n480,n479);
and gate_461(n481,n122,n461);
and gate_462(n482,n30,n481);
not gate_463(n483,n482);
and gate_464(n484,n480,n483);
not gate_465(n485,n484);
and gate_466(n486,n27,n485);
not gate_467(n487,n486);
and gate_468(n488,n476,n487);
not gate_469(n489,n488);
and gate_470(n490,n98,n489);
not gate_471(n491,n490);
and gate_472(n492,n460,n491);
and gate_473(n493,n387,n492);
not gate_474(n494,n493);
and gate_475(n495,n20,n494);
not gate_476(n496,n495);
and gate_477(n497,n349,n496);
not gate_478(n498,n497);
and gate_479(n499,n26,n498);
not gate_480(n500,n499);
and gate_481(n501,pi4,n188);
and gate_482(n502,n68,n501);
not gate_483(n503,n502);
and gate_484(n504,n24,n179);
not gate_485(n505,n504);
and gate_486(n506,pi4,n181);
not gate_487(n507,n506);
and gate_488(n508,n505,n507);
not gate_489(n509,n508);
and gate_490(n510,pi0,n337);
and gate_491(n511,n509,n510);
not gate_492(n512,n511);
and gate_493(n513,n503,n512);
not gate_494(n514,n513);
and gate_495(n515,n357,n514);
not gate_496(n516,n515);
and gate_497(n517,pi3,n278);
and gate_498(n518,n84,n517);
not gate_499(n519,n518);
and gate_500(n520,n20,n29);
not gate_501(n521,n520);
and gate_502(n522,n21,pi3);
not gate_503(n523,n522);
and gate_504(n524,n356,n523);
and gate_505(n525,n520,n524);
not gate_506(n526,n525);
and gate_507(n527,n519,n526);
not gate_508(n528,n527);
and gate_509(n529,n27,n528);
not gate_510(n530,n529);
and gate_511(n531,n20,pi3);
not gate_512(n532,n531);
and gate_513(n533,n39,n531);
not gate_514(n534,n533);
and gate_515(n535,pi0,pi9);
not gate_516(n536,n535);
and gate_517(n537,n521,n536);
not gate_518(n538,n537);
and gate_519(n539,n28,n537);
and gate_520(n540,n532,n539);
not gate_521(n541,n540);
and gate_522(n542,n534,n541);
not gate_523(n543,n542);
and gate_524(n544,pi1,pi7);
not gate_525(n545,n544);
and gate_526(n546,n543,n544);
not gate_527(n547,n546);
and gate_528(n548,n530,n547);
not gate_529(n549,n548);
and gate_530(n550,pi2,n549);
not gate_531(n551,n550);
and gate_532(n552,n21,pi7);
and gate_533(n553,n20,n552);
not gate_534(n554,n553);
and gate_535(n555,n233,n373);
not gate_536(n556,n555);
and gate_537(n557,pi0,n27);
not gate_538(n558,n557);
and gate_539(n559,n555,n558);
and gate_540(n560,n554,n559);
and gate_541(n561,pi9,n560);
not gate_542(n562,n561);
and gate_543(n563,n77,n85);
not gate_544(n564,n563);
and gate_545(n565,pi1,pi8);
not gate_546(n566,n565);
and gate_547(n567,n21,n28);
not gate_548(n568,n567);
and gate_549(n569,n566,n568);
not gate_550(n570,n569);
and gate_551(n571,n190,n570);
and gate_552(n572,n563,n571);
not gate_553(n573,n572);
and gate_554(n574,n562,n573);
not gate_555(n575,n574);
and gate_556(n576,pi3,n575);
not gate_557(n577,n576);
and gate_558(n578,pi1,pi9);
not gate_559(n579,n578);
and gate_560(n580,n21,n29);
not gate_561(n581,n580);
and gate_562(n582,n579,n581);
not gate_563(n583,n582);
and gate_564(n584,pi0,n583);
not gate_565(n585,n584);
and gate_566(n586,pi1,n29);
not gate_567(n587,n586);
and gate_568(n588,n20,n586);
not gate_569(n589,n588);
and gate_570(n590,n585,n589);
not gate_571(n591,n590);
and gate_572(n592,n23,n419);
and gate_573(n593,n591,n592);
not gate_574(n594,n593);
and gate_575(n595,n577,n594);
not gate_576(n596,n595);
and gate_577(n597,n22,n596);
not gate_578(n598,n597);
and gate_579(n599,n551,n598);
not gate_580(n600,n599);
and gate_581(n601,pi4,n600);
not gate_582(n602,n601);
and gate_583(n603,pi1,n285);
not gate_584(n604,n603);
and gate_585(n605,n21,n23);
and gate_586(n606,n39,n605);
not gate_587(n607,n606);
and gate_588(n608,n604,n607);
not gate_589(n609,n608);
and gate_590(n610,n22,n609);
not gate_591(n611,n610);
and gate_592(n612,pi2,n28);
not gate_593(n613,n612);
and gate_594(n614,n605,n612);
not gate_595(n615,n614);
and gate_596(n616,n611,n615);
not gate_597(n617,n616);
and gate_598(n618,pi7,n617);
not gate_599(n619,n618);
and gate_600(n620,pi3,pi9);
not gate_601(n621,n620);
and gate_602(n622,n27,n356);
and gate_603(n623,n621,n622);
and gate_604(n624,n104,n623);
not gate_605(n625,n624);
and gate_606(n626,n619,n625);
not gate_607(n627,n626);
and gate_608(n628,n20,n627);
not gate_609(n629,n628);
and gate_610(n630,n22,pi8);
not gate_611(n631,n630);
and gate_612(n632,n613,n631);
not gate_613(n633,n632);
and gate_614(n634,pi1,n633);
not gate_615(n635,n634);
and gate_616(n636,pi2,pi8);
not gate_617(n637,n636);
and gate_618(n638,n21,n636);
not gate_619(n639,n638);
and gate_620(n640,n635,n639);
not gate_621(n641,n640);
and gate_622(n642,pi3,n641);
not gate_623(n643,n642);
and gate_624(n644,pi1,n22);
not gate_625(n645,n644);
and gate_626(n646,n327,n644);
not gate_627(n647,n646);
and gate_628(n648,n643,n647);
not gate_629(n649,n648);
and gate_630(n650,n190,n649);
and gate_631(n651,pi0,n650);
not gate_632(n652,n651);
and gate_633(n653,n629,n652);
not gate_634(n654,n653);
and gate_635(n655,n24,n654);
not gate_636(n656,n655);
and gate_637(n657,n602,n656);
and gate_638(n658,n516,n657);
not gate_639(n659,n658);
and gate_640(n660,pi5,n659);
not gate_641(n661,n660);
and gate_642(n662,n20,pi2);
and gate_643(n663,n501,n662);
not gate_644(n664,n663);
and gate_645(n665,n82,n363);
and gate_646(n666,n114,n665);
not gate_647(n667,n666);
and gate_648(n668,n664,n667);
not gate_649(n669,n668);
and gate_650(n670,n330,n669);
not gate_651(n671,n670);
and gate_652(n672,n22,pi9);
not gate_653(n673,n672);
and gate_654(n674,pi0,n672);
not gate_655(n675,n674);
and gate_656(n676,pi2,n29);
not gate_657(n677,n676);
and gate_658(n678,n20,n676);
not gate_659(n679,n678);
and gate_660(n680,n675,n679);
not gate_661(n681,n680);
and gate_662(n682,n20,n380);
not gate_663(n683,n682);
and gate_664(n684,n680,n683);
not gate_665(n685,n684);
and gate_666(n686,n27,n685);
not gate_667(n687,n686);
and gate_668(n688,n24,pi7);
not gate_669(n689,n688);
and gate_670(n690,n20,n22);
not gate_671(n691,n690);
and gate_672(n692,n688,n690);
not gate_673(n693,n692);
and gate_674(n694,n687,n693);
not gate_675(n695,n694);
and gate_676(n696,n28,n695);
not gate_677(n697,n696);
and gate_678(n698,pi2,pi4);
and gate_679(n699,n20,n698);
and gate_680(n700,pi7,n278);
not gate_681(n701,n700);
and gate_682(n702,n699,n700);
not gate_683(n703,n702);
and gate_684(n704,n697,n703);
not gate_685(n705,n704);
and gate_686(n706,pi3,n705);
not gate_687(n707,n706);
and gate_688(n708,pi4,n39);
not gate_689(n709,n708);
and gate_690(n710,n20,n708);
not gate_691(n711,n710);
and gate_692(n712,pi0,pi2);
not gate_693(n713,n712);
and gate_694(n714,n24,n32);
not gate_695(n715,n714);
and gate_696(n716,n712,n714);
not gate_697(n717,n716);
and gate_698(n718,n711,n717);
not gate_699(n719,n718);
and gate_700(n720,n448,n719);
not gate_701(n721,n720);
and gate_702(n722,n707,n721);
and gate_703(n723,n671,n722);
not gate_704(n724,n723);
and gate_705(n725,n21,n724);
not gate_706(n726,n725);
and gate_707(n727,pi3,pi7);
not gate_708(n728,n727);
and gate_709(n729,n449,n728);
not gate_710(n730,n729);
and gate_711(n731,pi2,n730);
not gate_712(n732,n731);
and gate_713(n733,n22,n255);
not gate_714(n734,n733);
and gate_715(n735,n732,n734);
not gate_716(n736,n735);
and gate_717(n737,n29,n736);
not gate_718(n738,n737);
and gate_719(n739,n179,n288);
not gate_720(n740,n739);
and gate_721(n741,n738,n740);
not gate_722(n742,n741);
and gate_723(n743,n28,n742);
not gate_724(n744,n743);
and gate_725(n745,n288,n307);
not gate_726(n746,n745);
and gate_727(n747,n744,n746);
not gate_728(n748,n747);
and gate_729(n749,pi4,n748);
not gate_730(n750,n749);
and gate_731(n751,n279,n364);
not gate_732(n752,n751);
and gate_733(n753,n248,n289);
not gate_734(n754,n753);
and gate_735(n755,n752,n754);
and gate_736(n756,n688,n755);
not gate_737(n757,n756);
and gate_738(n758,n750,n757);
not gate_739(n759,n758);
and gate_740(n760,pi0,n759);
not gate_741(n761,n760);
and gate_742(n762,pi4,pi9);
not gate_743(n763,n762);
and gate_744(n764,pi3,n762);
not gate_745(n765,n764);
and gate_746(n766,n24,n29);
not gate_747(n767,n766);
and gate_748(n768,n23,n766);
not gate_749(n769,n768);
and gate_750(n770,n765,n769);
not gate_751(n771,n770);
and gate_752(n772,n22,n28);
not gate_753(n773,n772);
and gate_754(n774,n771,n772);
not gate_755(n775,n774);
and gate_756(n776,n23,n240);
not gate_757(n777,n776);
and gate_758(n778,pi8,n777);
and gate_759(n779,n80,n778);
not gate_760(n780,n779);
and gate_761(n781,n775,n780);
not gate_762(n782,n781);
and gate_763(n783,pi7,n782);
not gate_764(n784,n783);
and gate_765(n785,n23,pi4);
not gate_766(n786,n785);
and gate_767(n787,pi2,n785);
and gate_768(n788,n267,n787);
not gate_769(n789,n788);
and gate_770(n790,n784,n789);
not gate_771(n791,n790);
and gate_772(n792,n20,n791);
not gate_773(n793,n792);
and gate_774(n794,n761,n793);
not gate_775(n795,n794);
and gate_776(n796,pi1,n795);
not gate_777(n797,n796);
and gate_778(n798,n726,n797);
not gate_779(n799,n798);
and gate_780(n800,n25,n799);
not gate_781(n801,n800);
and gate_782(n802,n661,n801);
not gate_783(n803,n802);
and gate_784(n804,pi6,n803);
not gate_785(n805,n804);
and gate_786(n806,n500,n805);
and gate_787(n807,n178,n806);
and gate_788(n808,n65,n807);
not gate_789(po0,n808);
and gate_790(n810,n265,n305);
not gate_791(n811,n810);
and gate_792(n812,n31,n810);
and gate_793(n813,n363,n812);
and gate_794(n814,n29,n813);
not gate_795(n815,n814);
and gate_796(n816,pi2,n408);
not gate_797(n817,n816);
and gate_798(n818,n815,n817);
not gate_799(n819,n818);
and gate_800(n820,pi1,n819);
not gate_801(n821,n820);
and gate_802(n822,n25,pi9);
not gate_803(n823,n822);
and gate_804(n824,pi3,n822);
not gate_805(n825,n824);
and gate_806(n826,n23,n121);
not gate_807(n827,n826);
and gate_808(n828,n825,n827);
not gate_809(n829,n828);
and gate_810(n830,pi2,n829);
not gate_811(n831,n830);
and gate_812(n832,pi5,pi9);
not gate_813(n833,n832);
and gate_814(n834,n288,n832);
not gate_815(n835,n834);
and gate_816(n836,n831,n835);
not gate_817(n837,n836);
and gate_818(n838,pi7,n837);
not gate_819(n839,n838);
and gate_820(n840,pi3,pi5);
not gate_821(n841,n840);
and gate_822(n842,n23,n25);
not gate_823(n843,n842);
and gate_824(n844,n841,n843);
not gate_825(n845,n844);
and gate_826(n846,n22,n188);
not gate_827(n847,n846);
and gate_828(n848,n845,n846);
not gate_829(n849,n848);
and gate_830(n850,n839,n849);
not gate_831(n851,n850);
and gate_832(n852,n21,n851);
not gate_833(n853,n852);
and gate_834(n854,n821,n853);
not gate_835(n855,n854);
and gate_836(n856,n20,n855);
not gate_837(n857,n856);
and gate_838(n858,n174,n240);
not gate_839(n859,n858);
and gate_840(n860,pi1,n858);
not gate_841(n861,n860);
and gate_842(n862,n31,n338);
and gate_843(n863,n861,n862);
and gate_844(n864,n27,n863);
not gate_845(n865,n864);
and gate_846(n866,n66,n190);
not gate_847(n867,n866);
and gate_848(n868,pi3,n866);
not gate_849(n869,n868);
and gate_850(n870,n865,n869);
not gate_851(n871,n870);
and gate_852(n872,pi5,n871);
not gate_853(n873,n872);
and gate_854(n874,pi2,n23);
and gate_855(n875,n21,n874);
and gate_856(n876,n25,n179);
and gate_857(n877,n875,n876);
not gate_858(n878,n877);
and gate_859(n879,n873,n878);
not gate_860(n880,n879);
and gate_861(n881,pi0,n880);
not gate_862(n882,n881);
and gate_863(n883,n857,n882);
not gate_864(n884,n883);
and gate_865(n885,pi4,n884);
not gate_866(n886,n885);
and gate_867(n887,n21,n466);
not gate_868(n888,n887);
and gate_869(n889,n22,pi5);
not gate_870(n890,n889);
and gate_871(n891,pi1,n889);
not gate_872(n892,n891);
and gate_873(n893,n888,n892);
not gate_874(n894,n893);
and gate_875(n895,n27,n894);
not gate_876(n896,n895);
and gate_877(n897,pi1,n49);
not gate_878(n898,n897);
and gate_879(n899,n896,n898);
not gate_880(n900,n899);
and gate_881(n901,n29,n900);
not gate_882(n902,n901);
and gate_883(n903,pi2,n223);
not gate_884(n904,n903);
and gate_885(n905,n22,n56);
not gate_886(n906,n905);
and gate_887(n907,n904,n906);
not gate_888(n908,n907);
and gate_889(n909,n21,pi9);
not gate_890(n910,n909);
and gate_891(n911,n908,n909);
not gate_892(n912,n911);
and gate_893(n913,n902,n912);
not gate_894(n914,n913);
and gate_895(n915,n23,n914);
not gate_896(n916,n915);
and gate_897(n917,pi2,n25);
not gate_898(n918,n917);
and gate_899(n919,n890,n918);
not gate_900(n920,n919);
and gate_901(n921,pi9,n920);
and gate_902(n922,n21,n921);
not gate_903(n923,n922);
and gate_904(n924,n673,n677);
not gate_905(n925,n924);
and gate_906(n926,n122,n823);
not gate_907(n927,n926);
and gate_908(n928,pi1,n926);
and gate_909(n929,n925,n928);
not gate_910(n930,n929);
and gate_911(n931,n923,n930);
not gate_912(n932,n931);
and gate_913(n933,n27,n932);
not gate_914(n934,n933);
and gate_915(n935,n321,n644);
not gate_916(n936,n935);
and gate_917(n937,n934,n936);
not gate_918(n938,n937);
and gate_919(n939,pi3,n938);
not gate_920(n940,n939);
and gate_921(n941,n916,n940);
not gate_922(n942,n941);
and gate_923(n943,n20,n942);
not gate_924(n944,n943);
and gate_925(n945,pi1,n23);
not gate_926(n946,n945);
and gate_927(n947,n832,n945);
not gate_928(n948,n947);
and gate_929(n949,n25,n29);
not gate_930(n950,n949);
and gate_931(n951,n833,n950);
not gate_932(n952,n951);
and gate_933(n953,n21,n858);
and gate_934(n954,n952,n953);
not gate_935(n955,n954);
and gate_936(n956,n948,n955);
not gate_937(n957,n956);
and gate_938(n958,n22,n957);
not gate_939(n959,n958);
and gate_940(n960,n23,n29);
not gate_941(n961,n960);
and gate_942(n962,n621,n961);
not gate_943(n963,n962);
and gate_944(n964,n917,n963);
and gate_945(n965,pi1,n964);
not gate_946(n966,n965);
and gate_947(n967,n959,n966);
not gate_948(n968,n967);
and gate_949(n969,n557,n968);
not gate_950(n970,n969);
and gate_951(n971,n944,n970);
not gate_952(n972,n971);
and gate_953(n973,n24,n972);
not gate_954(n974,n973);
and gate_955(n975,n886,n974);
not gate_956(n976,n975);
and gate_957(n977,n26,n976);
not gate_958(n978,n977);
and gate_959(n979,pi4,pi5);
not gate_960(n980,n979);
and gate_961(n981,n522,n979);
not gate_962(n982,n981);
and gate_963(n983,n24,n25);
not gate_964(n984,n983);
and gate_965(n985,n945,n983);
not gate_966(n986,n985);
and gate_967(n987,n982,n986);
not gate_968(n988,n987);
and gate_969(n989,n691,n713);
not gate_970(n990,n989);
and gate_971(n991,n988,n990);
not gate_972(n992,n991);
and gate_973(n993,n21,n785);
not gate_974(n994,n993);
and gate_975(n995,pi3,n24);
not gate_976(n996,n995);
and gate_977(n997,pi1,n995);
not gate_978(n998,n997);
and gate_979(n999,n994,n998);
not gate_980(n1000,n999);
and gate_981(n1001,pi0,n1000);
not gate_982(n1002,n1001);
and gate_983(n1003,pi1,pi4);
not gate_984(n1004,n1003);
and gate_985(n1005,n21,n24);
not gate_986(n1006,n1005);
and gate_987(n1007,n1004,n1006);
not gate_988(n1008,n1007);
and gate_989(n1009,n531,n1008);
not gate_990(n1010,n1009);
and gate_991(n1011,n1002,n1010);
not gate_992(n1012,n1011);
and gate_993(n1013,n463,n1012);
not gate_994(n1014,n1013);
and gate_995(n1015,n992,n1014);
not gate_996(n1016,n1015);
and gate_997(n1017,pi9,n1016);
not gate_998(n1018,n1017);
and gate_999(n1019,n24,pi5);
not gate_1000(n1020,n1019);
and gate_1001(n1021,pi4,n25);
not gate_1002(n1022,n1021);
and gate_1003(n1023,n1020,n1022);
not gate_1004(n1024,n1023);
and gate_1005(n1025,pi1,n810);
and gate_1006(n1026,n1024,n1025);
not gate_1007(n1027,n1026);
and gate_1008(n1028,n982,n1027);
not gate_1009(n1029,n1028);
and gate_1010(n1030,n22,n1029);
not gate_1011(n1031,n1030);
and gate_1012(n1032,n104,n1019);
not gate_1013(n1033,n1032);
and gate_1014(n1034,n1031,n1033);
not gate_1015(n1035,n1034);
and gate_1016(n1036,pi0,n1035);
not gate_1017(n1037,n1036);
and gate_1018(n1038,n605,n983);
not gate_1019(n1039,n1038);
and gate_1020(n1040,n370,n980);
not gate_1021(n1041,n1040);
and gate_1022(n1042,pi3,n351);
and gate_1023(n1043,n1041,n1042);
not gate_1024(n1044,n1043);
and gate_1025(n1045,n1039,n1044);
not gate_1026(n1046,n1045);
and gate_1027(n1047,n662,n1046);
not gate_1028(n1048,n1047);
and gate_1029(n1049,n1037,n1048);
not gate_1030(n1050,n1049);
and gate_1031(n1051,n29,n1050);
not gate_1032(n1052,n1051);
and gate_1033(n1053,n1018,n1052);
not gate_1034(n1054,n1053);
and gate_1035(n1055,n27,n1054);
not gate_1036(n1056,n1055);
and gate_1037(n1057,n980,n984);
not gate_1038(n1058,n1057);
and gate_1039(n1059,n465,n1057);
and gate_1040(n1060,n351,n1059);
and gate_1041(n1061,n23,n1060);
not gate_1042(n1062,n1061);
and gate_1043(n1063,n21,n1021);
and gate_1044(n1064,n288,n1063);
not gate_1045(n1065,n1064);
and gate_1046(n1066,n1062,n1065);
not gate_1047(n1067,n1066);
and gate_1048(n1068,n20,n1067);
not gate_1049(n1069,n1068);
and gate_1050(n1070,pi0,n104);
and gate_1051(n1071,n786,n996);
not gate_1052(n1072,n1071);
and gate_1053(n1073,n984,n1071);
and gate_1054(n1074,n1070,n1073);
not gate_1055(n1075,n1074);
and gate_1056(n1076,n1069,n1075);
not gate_1057(n1077,n1076);
and gate_1058(n1078,n29,n1077);
not gate_1059(n1079,n1078);
and gate_1060(n1080,n690,n840);
not gate_1061(n1081,n1080);
and gate_1062(n1082,pi0,n919);
and gate_1063(n1083,n811,n1082);
not gate_1064(n1084,n1083);
and gate_1065(n1085,n1081,n1084);
not gate_1066(n1086,n1085);
and gate_1067(n1087,pi1,n1086);
not gate_1068(n1088,n1087);
and gate_1069(n1089,pi2,n264);
and gate_1070(n1090,n47,n1089);
not gate_1071(n1091,n1090);
and gate_1072(n1092,n1088,n1091);
not gate_1073(n1093,n1092);
and gate_1074(n1094,n24,n1093);
not gate_1075(n1095,n1094);
and gate_1076(n1096,n23,n1021);
and gate_1077(n1097,pi0,n66);
not gate_1078(n1098,n1097);
and gate_1079(n1099,n1096,n1097);
not gate_1080(n1100,n1099);
and gate_1081(n1101,n1095,n1100);
not gate_1082(n1102,n1101);
and gate_1083(n1103,pi9,n1102);
not gate_1084(n1104,n1103);
and gate_1085(n1105,n1079,n1104);
not gate_1086(n1106,n1105);
and gate_1087(n1107,pi7,n1106);
not gate_1088(n1108,n1107);
and gate_1089(n1109,n1056,n1108);
not gate_1090(n1110,n1109);
and gate_1091(n1111,pi6,n1110);
not gate_1092(n1112,n1111);
and gate_1093(n1113,n978,n1112);
and gate_1094(n1114,n105,n645);
not gate_1095(n1115,n1114);
and gate_1096(n1116,n58,n1115);
and gate_1097(n1117,n20,n1116);
not gate_1098(n1118,n1117);
and gate_1099(n1119,n51,n510);
not gate_1100(n1120,n1119);
and gate_1101(n1121,n1118,n1120);
not gate_1102(n1122,n1121);
and gate_1103(n1123,pi6,n29);
not gate_1104(n1124,n1123);
and gate_1105(n1125,n26,pi9);
not gate_1106(n1126,n1125);
and gate_1107(n1127,n1124,n1126);
not gate_1108(n1128,n1127);
and gate_1109(n1129,n1122,n1127);
and gate_1110(n1130,n859,n1129);
not gate_1111(n1131,n1130);
and gate_1112(n1132,n1113,n1131);
not gate_1113(n1133,n1132);
and gate_1114(n1134,n28,n1133);
not gate_1115(n1135,n1134);
and gate_1116(n1136,pi1,n83);
not gate_1117(n1137,n1136);
and gate_1118(n1138,n21,n698);
not gate_1119(n1139,n1138);
and gate_1120(n1140,n1137,n1139);
not gate_1121(n1141,n1140);
and gate_1122(n1142,pi6,n1141);
not gate_1123(n1143,n1142);
and gate_1124(n1144,n21,n26);
not gate_1125(n1145,n1144);
and gate_1126(n1146,n82,n1144);
not gate_1127(n1147,n1146);
and gate_1128(n1148,n1143,n1147);
not gate_1129(n1149,n1148);
and gate_1130(n1150,n29,n1149);
not gate_1131(n1151,n1150);
and gate_1132(n1152,pi4,pi6);
not gate_1133(n1153,n1152);
and gate_1134(n1154,n24,n26);
not gate_1135(n1155,n1154);
and gate_1136(n1156,n1153,n1155);
not gate_1137(n1157,n1156);
and gate_1138(n1158,n21,n1157);
not gate_1139(n1159,n1158);
and gate_1140(n1160,pi1,n106);
not gate_1141(n1161,n1160);
and gate_1142(n1162,n1159,n1161);
not gate_1143(n1163,n1162);
and gate_1144(n1164,pi2,pi9);
not gate_1145(n1165,n1164);
and gate_1146(n1166,n1163,n1164);
not gate_1147(n1167,n1166);
and gate_1148(n1168,n1151,n1167);
not gate_1149(n1169,n1168);
and gate_1150(n1170,pi7,n1169);
not gate_1151(n1171,n1170);
and gate_1152(n1172,n66,n380);
not gate_1153(n1173,n1172);
and gate_1154(n1174,n22,n29);
not gate_1155(n1175,n1174);
and gate_1156(n1176,n1165,n1175);
not gate_1157(n1177,n1176);
and gate_1158(n1178,n21,pi4);
not gate_1159(n1179,n1178);
and gate_1160(n1180,n1177,n1178);
not gate_1161(n1181,n1180);
and gate_1162(n1182,n1173,n1181);
not gate_1163(n1183,n1182);
and gate_1164(n1184,n26,n1183);
not gate_1165(n1185,n1184);
and gate_1166(n1186,n24,n1123);
and gate_1167(n1187,n337,n1186);
not gate_1168(n1188,n1187);
and gate_1169(n1189,n1185,n1188);
not gate_1170(n1190,n1189);
and gate_1171(n1191,n27,n1190);
not gate_1172(n1192,n1191);
and gate_1173(n1193,n1171,n1192);
not gate_1174(n1194,n1193);
and gate_1175(n1195,pi5,n1194);
not gate_1176(n1196,n1195);
and gate_1177(n1197,n26,pi7);
not gate_1178(n1198,n1197);
and gate_1179(n1199,n167,n1198);
not gate_1180(n1200,n1199);
and gate_1181(n1201,n67,n338);
not gate_1182(n1202,n1201);
and gate_1183(n1203,n1200,n1202);
and gate_1184(n1204,n24,n1203);
not gate_1185(n1205,n1204);
and gate_1186(n1206,pi4,n166);
not gate_1187(n1207,n1206);
and gate_1188(n1208,n21,n1206);
not gate_1189(n1209,n1208);
and gate_1190(n1210,n1205,n1209);
not gate_1191(n1211,n1210);
and gate_1192(n1212,n29,n1211);
not gate_1193(n1213,n1212);
and gate_1194(n1214,n21,pi6);
not gate_1195(n1215,n1214);
and gate_1196(n1216,n188,n1214);
not gate_1197(n1217,n1216);
and gate_1198(n1218,n80,n1216);
not gate_1199(n1219,n1218);
and gate_1200(n1220,n1213,n1219);
not gate_1201(n1221,n1220);
and gate_1202(n1222,n25,n1221);
not gate_1203(n1223,n1222);
and gate_1204(n1224,n1196,n1223);
not gate_1205(n1225,n1224);
and gate_1206(n1226,pi0,n1225);
not gate_1207(n1227,n1226);
and gate_1208(n1228,n1137,n1215);
not gate_1209(n1229,n1228);
and gate_1210(n1230,n1156,n1229);
and gate_1211(n1231,pi9,n1230);
not gate_1212(n1232,n1231);
and gate_1213(n1233,n24,pi6);
not gate_1214(n1234,n1233);
and gate_1215(n1235,n107,n1234);
not gate_1216(n1236,n1235);
and gate_1217(n1237,n81,n1235);
and gate_1218(n1238,n580,n1237);
not gate_1219(n1239,n1238);
and gate_1220(n1240,n1232,n1239);
not gate_1221(n1241,n1240);
and gate_1222(n1242,n25,n1241);
not gate_1223(n1243,n1242);
and gate_1224(n1244,pi1,n123);
not gate_1225(n1245,n1244);
and gate_1226(n1246,n21,n124);
not gate_1227(n1247,n1246);
and gate_1228(n1248,n1245,n1247);
and gate_1229(n1249,n1156,n1248);
and gate_1230(n1250,n889,n1249);
not gate_1231(n1251,n1250);
and gate_1232(n1252,n1243,n1251);
not gate_1233(n1253,n1252);
and gate_1234(n1254,pi7,n1253);
not gate_1235(n1255,n1254);
and gate_1236(n1256,n644,n1236);
not gate_1237(n1257,n1256);
and gate_1238(n1258,n109,n1257);
not gate_1239(n1259,n1258);
and gate_1240(n1260,pi9,n1259);
not gate_1241(n1261,n1260);
and gate_1242(n1262,n104,n1186);
not gate_1243(n1263,n1262);
and gate_1244(n1264,n1261,n1263);
not gate_1245(n1265,n1264);
and gate_1246(n1266,n153,n1265);
not gate_1247(n1267,n1266);
and gate_1248(n1268,n1255,n1267);
not gate_1249(n1269,n1268);
and gate_1250(n1270,n20,n1269);
not gate_1251(n1271,n1270);
and gate_1252(n1272,n1227,n1271);
not gate_1253(n1273,n1272);
and gate_1254(n1274,n23,n1273);
not gate_1255(n1275,n1274);
and gate_1256(n1276,n25,n1125);
and gate_1257(n1277,n644,n1276);
not gate_1258(n1278,n1277);
and gate_1259(n1279,pi5,n1123);
and gate_1260(n1280,n104,n1279);
not gate_1261(n1281,n1280);
and gate_1262(n1282,n1278,n1281);
not gate_1263(n1283,n1282);
and gate_1264(n1284,n24,n1283);
and gate_1265(n1285,pi0,n1284);
not gate_1266(n1286,n1285);
and gate_1267(n1287,n20,n337);
and gate_1268(n1288,n979,n1123);
and gate_1269(n1289,n1287,n1288);
not gate_1270(n1290,n1289);
and gate_1271(n1291,n1286,n1290);
and gate_1272(n1292,n20,pi4);
and gate_1273(n1293,n26,n179);
not gate_1274(n1294,n1293);
and gate_1275(n1295,n1292,n1293);
not gate_1276(n1296,n1295);
and gate_1277(n1297,n20,pi7);
not gate_1278(n1298,n1297);
and gate_1279(n1299,n558,n1298);
not gate_1280(n1300,n1299);
and gate_1281(n1301,n1236,n1300);
and gate_1282(n1302,n193,n1301);
not gate_1283(n1303,n1302);
and gate_1284(n1304,n1296,n1303);
not gate_1285(n1305,n1304);
and gate_1286(n1306,pi1,n1305);
not gate_1287(n1307,n1306);
and gate_1288(n1308,pi0,pi6);
not gate_1289(n1309,n1308);
and gate_1290(n1310,n189,n1299);
and gate_1291(n1311,n1309,n1310);
and gate_1292(n1312,n1178,n1311);
not gate_1293(n1313,n1312);
and gate_1294(n1314,n1307,n1313);
not gate_1295(n1315,n1314);
and gate_1296(n1316,pi5,n1315);
not gate_1297(n1317,n1316);
and gate_1298(n1318,pi4,n822);
not gate_1299(n1319,n1318);
and gate_1300(n1320,pi6,pi7);
not gate_1301(n1321,n1320);
and gate_1302(n1322,n21,n1320);
not gate_1303(n1323,n1322);
and gate_1304(n1324,n26,n27);
not gate_1305(n1325,n1324);
and gate_1306(n1326,pi1,n1324);
not gate_1307(n1327,n1326);
and gate_1308(n1328,n1323,n1327);
not gate_1309(n1329,n1328);
and gate_1310(n1330,pi0,n1329);
not gate_1311(n1331,n1330);
and gate_1312(n1332,pi1,n26);
not gate_1313(n1333,n1332);
and gate_1314(n1334,n1215,n1333);
not gate_1315(n1335,n1334);
and gate_1316(n1336,n20,n27);
not gate_1317(n1337,n1336);
and gate_1318(n1338,n1334,n1336);
not gate_1319(n1339,n1338);
and gate_1320(n1340,n1331,n1339);
not gate_1321(n1341,n1340);
and gate_1322(n1342,n1318,n1341);
not gate_1323(n1343,n1342);
and gate_1324(n1344,n1317,n1343);
not gate_1325(n1345,n1344);
and gate_1326(n1346,pi2,n1345);
not gate_1327(n1347,n1346);
and gate_1328(n1348,n27,n1236);
and gate_1329(n1349,n1334,n1348);
and gate_1330(n1350,pi0,n1349);
not gate_1331(n1351,n1350);
and gate_1332(n1352,n21,n1197);
and gate_1333(n1353,n20,n1352);
not gate_1334(n1354,n1353);
and gate_1335(n1355,n1351,n1354);
not gate_1336(n1356,n1355);
and gate_1337(n1357,pi9,n1356);
not gate_1338(n1358,n1357);
and gate_1339(n1359,pi0,n98);
and gate_1340(n1360,pi6,n181);
not gate_1341(n1361,n1360);
and gate_1342(n1362,n1359,n1360);
not gate_1343(n1363,n1362);
and gate_1344(n1364,n1358,n1363);
not gate_1345(n1365,n1364);
and gate_1346(n1366,n889,n1365);
not gate_1347(n1367,n1366);
and gate_1348(n1368,n1347,n1367);
and gate_1349(n1369,n74,n1276);
not gate_1350(n1370,n1369);
and gate_1351(n1371,n80,n1279);
not gate_1352(n1372,n1371);
and gate_1353(n1373,n1370,n1372);
not gate_1354(n1374,n1373);
and gate_1355(n1375,n563,n1374);
and gate_1356(n1376,n1300,n1375);
not gate_1357(n1377,n1376);
and gate_1358(n1378,n1368,n1377);
and gate_1359(n1379,n1291,n1378);
not gate_1360(n1380,n1379);
and gate_1361(n1381,pi3,n1380);
not gate_1362(n1382,n1381);
and gate_1363(n1383,n1275,n1382);
not gate_1364(n1384,n1383);
and gate_1365(n1385,pi8,n1384);
not gate_1366(n1386,n1385);
and gate_1367(n1387,n1135,n1386);
not gate_1368(po1,n1387);
and gate_1369(n1389,pi3,n99);
and gate_1370(n1390,n104,n1389);
not gate_1371(n1391,n1390);
and gate_1372(n1392,n70,n91);
not gate_1373(n1393,n1392);
and gate_1374(n1394,n466,n1393);
and gate_1375(n1395,n945,n1394);
not gate_1376(n1396,n1395);
and gate_1377(n1397,n1391,n1396);
not gate_1378(n1398,n1397);
and gate_1379(n1399,n509,n1398);
not gate_1380(n1400,n1399);
and gate_1381(n1401,n1294,n1361);
not gate_1382(n1402,n1401);
and gate_1383(n1403,n21,n1402);
not gate_1384(n1404,n1403);
and gate_1385(n1405,n181,n1332);
not gate_1386(n1406,n1405);
and gate_1387(n1407,n1404,n1406);
not gate_1388(n1408,n1407);
and gate_1389(n1409,pi4,n1408);
not gate_1390(n1410,n1409);
and gate_1391(n1411,n189,n1321);
not gate_1392(n1412,n1411);
and gate_1393(n1413,n98,n1412);
not gate_1394(n1414,n1413);
and gate_1395(n1415,n1410,n1414);
not gate_1396(n1416,n1415);
and gate_1397(n1417,pi2,n1416);
not gate_1398(n1418,n1417);
and gate_1399(n1419,pi1,pi6);
not gate_1400(n1420,n1419);
and gate_1401(n1421,pi4,n27);
not gate_1402(n1422,n1421);
and gate_1403(n1423,n689,n1422);
not gate_1404(n1424,n1423);
and gate_1405(n1425,n384,n1424);
and gate_1406(n1426,n1419,n1425);
not gate_1407(n1427,n1426);
and gate_1408(n1428,n21,n1324);
not gate_1409(n1429,n1428);
and gate_1410(n1430,n383,n1428);
not gate_1411(n1431,n1430);
and gate_1412(n1432,n1427,n1431);
not gate_1413(n1433,n1432);
and gate_1414(n1434,n22,n1433);
not gate_1415(n1435,n1434);
and gate_1416(n1436,n1418,n1435);
not gate_1417(n1437,n1436);
and gate_1418(n1438,n23,n1437);
not gate_1419(n1439,n1438);
and gate_1420(n1440,n21,n358);
not gate_1421(n1441,n1440);
and gate_1422(n1442,pi2,pi6);
not gate_1423(n1443,n1442);
and gate_1424(n1444,pi1,n1443);
and gate_1425(n1445,n359,n1198);
and gate_1426(n1446,n1444,n1445);
not gate_1427(n1447,n1446);
and gate_1428(n1448,n1441,n1447);
not gate_1429(n1449,n1448);
and gate_1430(n1450,n24,n1449);
not gate_1431(n1451,n1450);
and gate_1432(n1452,n1321,n1325);
not gate_1433(n1453,n1452);
and gate_1434(n1454,pi2,n1453);
not gate_1435(n1455,n1454);
and gate_1436(n1456,n1003,n1454);
not gate_1437(n1457,n1456);
and gate_1438(n1458,n1451,n1457);
not gate_1439(n1459,n1458);
and gate_1440(n1460,n29,n1459);
not gate_1441(n1461,n1460);
and gate_1442(n1462,n337,n1320);
not gate_1443(n1463,n1462);
and gate_1444(n1464,n1447,n1463);
not gate_1445(n1465,n1464);
and gate_1446(n1466,n762,n1465);
not gate_1447(n1467,n1466);
and gate_1448(n1468,n1461,n1467);
not gate_1449(n1469,n1468);
and gate_1450(n1470,pi3,n1469);
not gate_1451(n1471,n1470);
and gate_1452(n1472,n1439,n1471);
not gate_1453(n1473,n1472);
and gate_1454(n1474,n25,n1473);
not gate_1455(n1475,n1474);
and gate_1456(n1476,pi1,pi3);
not gate_1457(n1477,n1476);
and gate_1458(n1478,n179,n1476);
not gate_1459(n1479,n1478);
and gate_1460(n1480,n21,n27);
not gate_1461(n1481,n1480);
and gate_1462(n1482,n545,n1481);
not gate_1463(n1483,n1482);
and gate_1464(n1484,n859,n1483);
and gate_1465(n1485,n26,n1484);
not gate_1466(n1486,n1485);
and gate_1467(n1487,n1479,n1486);
not gate_1468(n1488,n1487);
and gate_1469(n1489,n22,n1488);
not gate_1470(n1490,n1489);
and gate_1471(n1491,pi3,n27);
not gate_1472(n1492,n1491);
and gate_1473(n1493,n21,n179);
not gate_1474(n1494,n1493);
and gate_1475(n1495,n1492,n1494);
not gate_1476(n1496,n1495);
and gate_1477(n1497,n523,n1496);
and gate_1478(n1498,n1442,n1497);
not gate_1479(n1499,n1498);
and gate_1480(n1500,n1490,n1499);
not gate_1481(n1501,n1500);
and gate_1482(n1502,n24,n1501);
not gate_1483(n1503,n1502);
and gate_1484(n1504,pi3,pi6);
not gate_1485(n1505,n1504);
and gate_1486(n1506,n23,n26);
not gate_1487(n1507,n1506);
and gate_1488(n1508,n1505,n1507);
not gate_1489(n1509,n1508);
and gate_1490(n1510,n22,n26);
not gate_1491(n1511,n1510);
and gate_1492(n1512,n1443,n1511);
not gate_1493(n1513,n1512);
and gate_1494(n1514,n1508,n1512);
and gate_1495(n1515,n1453,n1514);
and gate_1496(n1516,pi1,n1515);
not gate_1497(n1517,n1516);
and gate_1498(n1518,n166,n874);
not gate_1499(n1519,n1518);
and gate_1500(n1520,n730,n1510);
not gate_1501(n1521,n1520);
and gate_1502(n1522,n1519,n1521);
not gate_1503(n1523,n1522);
and gate_1504(n1524,n21,n1523);
not gate_1505(n1525,n1524);
and gate_1506(n1526,n1517,n1525);
not gate_1507(n1527,n1526);
and gate_1508(n1528,pi9,n1527);
not gate_1509(n1529,n1528);
and gate_1510(n1530,n23,n190);
and gate_1511(n1531,n1214,n1530);
not gate_1512(n1532,n1531);
and gate_1513(n1533,n1529,n1532);
not gate_1514(n1534,n1533);
and gate_1515(n1535,pi4,n1534);
not gate_1516(n1536,n1535);
and gate_1517(n1537,n1503,n1536);
not gate_1518(n1538,n1537);
and gate_1519(n1539,pi5,n1538);
not gate_1520(n1540,n1539);
and gate_1521(n1541,n1475,n1540);
and gate_1522(n1542,n1400,n1541);
not gate_1523(n1543,n1542);
and gate_1524(n1544,n28,n1543);
not gate_1525(n1545,n1544);
and gate_1526(n1546,n188,n337);
not gate_1527(n1547,n1546);
and gate_1528(n1548,n867,n1547);
not gate_1529(n1549,n1548);
and gate_1530(n1550,n1393,n1549);
not gate_1531(n1551,n1550);
and gate_1532(n1552,pi6,n190);
and gate_1533(n1553,n21,n917);
not gate_1534(n1554,n1553);
and gate_1535(n1555,n1552,n1553);
not gate_1536(n1556,n1555);
and gate_1537(n1557,n22,n1200);
not gate_1538(n1558,n1557);
and gate_1539(n1559,n1455,n1558);
not gate_1540(n1560,n1559);
and gate_1541(n1561,n25,n1560);
not gate_1542(n1562,n1561);
and gate_1543(n1563,n889,n1197);
not gate_1544(n1564,n1563);
and gate_1545(n1565,n1562,n1564);
not gate_1546(n1566,n1565);
and gate_1547(n1567,n578,n1566);
not gate_1548(n1568,n1567);
and gate_1549(n1569,n1556,n1568);
and gate_1550(n1570,n1551,n1569);
not gate_1551(n1571,n1570);
and gate_1552(n1572,n24,n1571);
not gate_1553(n1573,n1572);
and gate_1554(n1574,n22,n1452);
not gate_1555(n1575,n1574);
and gate_1556(n1576,n91,n918);
and gate_1557(n1577,n1575,n1576);
and gate_1558(n1578,pi9,n1577);
not gate_1559(n1579,n1578);
and gate_1560(n1580,n463,n1552);
not gate_1561(n1581,n1580);
and gate_1562(n1582,n1579,n1581);
not gate_1563(n1583,n1582);
and gate_1564(n1584,n21,n1583);
not gate_1565(n1585,n1584);
and gate_1566(n1586,pi6,n179);
not gate_1567(n1587,n1586);
and gate_1568(n1588,pi1,n463);
and gate_1569(n1589,n1586,n1588);
not gate_1570(n1590,n1589);
and gate_1571(n1591,n1585,n1590);
not gate_1572(n1592,n1591);
and gate_1573(n1593,pi4,n1592);
not gate_1574(n1594,n1593);
and gate_1575(n1595,n1573,n1594);
not gate_1576(n1596,n1595);
and gate_1577(n1597,pi3,n1596);
not gate_1578(n1598,n1597);
and gate_1579(n1599,pi5,n190);
and gate_1580(n1600,n24,n1599);
not gate_1581(n1601,n1600);
and gate_1582(n1602,pi9,n689);
and gate_1583(n1603,n980,n1602);
not gate_1584(n1604,n1603);
and gate_1585(n1605,n1601,n1604);
not gate_1586(n1606,n1605);
and gate_1587(n1607,n26,n1606);
not gate_1588(n1608,n1607);
and gate_1589(n1609,pi5,n1320);
and gate_1590(n1610,n381,n1609);
not gate_1591(n1611,n1610);
and gate_1592(n1612,n1608,n1611);
not gate_1593(n1613,n1612);
and gate_1594(n1614,pi2,n1613);
not gate_1595(n1615,n1614);
and gate_1596(n1616,n22,n979);
and gate_1597(n1617,n1293,n1616);
not gate_1598(n1618,n1617);
and gate_1599(n1619,n1615,n1618);
not gate_1600(n1620,n1619);
and gate_1601(n1621,pi1,n1620);
not gate_1602(n1622,n1621);
and gate_1603(n1623,pi2,n1153);
not gate_1604(n1624,n1623);
and gate_1605(n1625,pi5,n26);
not gate_1606(n1626,n1625);
and gate_1607(n1627,n100,n1626);
not gate_1608(n1628,n1627);
and gate_1609(n1629,n1155,n1627);
and gate_1610(n1630,n1624,n1629);
and gate_1611(n1631,n188,n1630);
and gate_1612(n1632,n21,n1631);
not gate_1613(n1633,n1632);
and gate_1614(n1634,n1622,n1633);
not gate_1615(n1635,n1634);
and gate_1616(n1636,n23,n1635);
not gate_1617(n1637,n1636);
and gate_1618(n1638,n1598,n1637);
and gate_1619(n1639,pi3,n1125);
not gate_1620(n1640,n1639);
and gate_1621(n1641,n23,n1123);
not gate_1622(n1642,n1641);
and gate_1623(n1643,n1640,n1642);
not gate_1624(n1644,n1643);
and gate_1625(n1645,n1021,n1644);
and gate_1626(n1646,pi2,n1645);
not gate_1627(n1647,n1646);
and gate_1628(n1648,n22,n995);
not gate_1629(n1649,n1648);
and gate_1630(n1650,pi5,n133);
and gate_1631(n1651,n1648,n1650);
not gate_1632(n1652,n1651);
and gate_1633(n1653,n1647,n1652);
not gate_1634(n1654,n1653);
and gate_1635(n1655,n1482,n1654);
not gate_1636(n1656,n1655);
and gate_1637(n1657,n1638,n1656);
not gate_1638(n1658,n1657);
and gate_1639(n1659,pi8,n1658);
not gate_1640(n1660,n1659);
and gate_1641(n1661,n1545,n1660);
not gate_1642(n1662,n1661);
and gate_1643(n1663,pi0,n1662);
not gate_1644(n1664,n1663);
and gate_1645(n1665,n23,n24);
not gate_1646(n1666,n1665);
and gate_1647(n1667,n21,n1665);
and gate_1648(n1668,n26,n28);
not gate_1649(n1669,n1668);
and gate_1650(n1670,pi5,n1668);
not gate_1651(n1671,n1670);
and gate_1652(n1672,n1667,n1670);
not gate_1653(n1673,n1672);
and gate_1654(n1674,pi6,pi8);
not gate_1655(n1675,n1674);
and gate_1656(n1676,n25,n1674);
not gate_1657(n1677,n1676);
and gate_1658(n1678,n1476,n1676);
not gate_1659(n1679,n1678);
and gate_1660(n1680,pi4,n1678);
not gate_1661(n1681,n1680);
and gate_1662(n1682,n1673,n1681);
not gate_1663(n1683,n1682);
and gate_1664(n1684,n29,n1683);
not gate_1665(n1685,n1684);
and gate_1666(n1686,n24,pi8);
not gate_1667(n1687,n1686);
and gate_1668(n1688,n522,n1686);
not gate_1669(n1689,n1688);
and gate_1670(n1690,pi4,n28);
not gate_1671(n1691,n1690);
and gate_1672(n1692,n945,n1690);
not gate_1673(n1693,n1692);
and gate_1674(n1694,n1689,n1693);
and gate_1675(n1695,n26,pi8);
not gate_1676(n1696,n1695);
and gate_1677(n1697,n23,n1695);
and gate_1678(n1698,n1003,n1697);
not gate_1679(n1699,n1698);
and gate_1680(n1700,n1694,n1699);
not gate_1681(n1701,n1700);
and gate_1682(n1702,pi5,n1701);
not gate_1683(n1703,n1702);
and gate_1684(n1704,pi4,pi8);
not gate_1685(n1705,n1704);
and gate_1686(n1706,n24,n28);
not gate_1687(n1707,n1706);
and gate_1688(n1708,n1705,n1707);
not gate_1689(n1709,n1708);
and gate_1690(n1710,pi1,n1709);
not gate_1691(n1711,n1710);
and gate_1692(n1712,n1006,n1711);
not gate_1693(n1713,n1712);
and gate_1694(n1714,n23,n69);
not gate_1695(n1715,n1714);
and gate_1696(n1716,n1713,n1714);
not gate_1697(n1717,n1716);
and gate_1698(n1718,n1703,n1717);
not gate_1699(n1719,n1718);
and gate_1700(n1720,pi9,n1719);
not gate_1701(n1721,n1720);
and gate_1702(n1722,n1685,n1721);
not gate_1703(n1723,n1722);
and gate_1704(n1724,pi2,n1723);
not gate_1705(n1725,n1724);
and gate_1706(n1726,n845,n1668);
and gate_1707(n1727,n21,n1726);
not gate_1708(n1728,n1727);
and gate_1709(n1729,n1679,n1728);
not gate_1710(n1730,n1729);
and gate_1711(n1731,n763,n767);
not gate_1712(n1732,n1731);
and gate_1713(n1733,n1730,n1732);
not gate_1714(n1734,n1733);
and gate_1715(n1735,n41,n842);
not gate_1716(n1736,n1735);
and gate_1717(n1737,pi6,n28);
not gate_1718(n1738,n1737);
and gate_1719(n1739,n1696,n1738);
not gate_1720(n1740,n1739);
and gate_1721(n1741,pi9,n1740);
and gate_1722(n1742,n811,n1741);
not gate_1723(n1743,n1742);
and gate_1724(n1744,n1736,n1743);
not gate_1725(n1745,n1744);
and gate_1726(n1746,pi4,n1745);
not gate_1727(n1747,n1746);
and gate_1728(n1748,n1669,n1675);
not gate_1729(n1749,n1748);
and gate_1730(n1750,n24,n121);
not gate_1731(n1751,n1750);
and gate_1732(n1752,n1749,n1750);
and gate_1733(n1753,n23,n1752);
not gate_1734(n1754,n1753);
and gate_1735(n1755,n1747,n1754);
not gate_1736(n1756,n1755);
and gate_1737(n1757,pi1,n1756);
not gate_1738(n1758,n1757);
and gate_1739(n1759,pi9,n330);
and gate_1740(n1760,n810,n1759);
and gate_1741(n1761,n1214,n1760);
not gate_1742(n1762,n1761);
and gate_1743(n1763,n1758,n1762);
and gate_1744(n1764,n1734,n1763);
not gate_1745(n1765,n1764);
and gate_1746(n1766,n22,n1765);
not gate_1747(n1767,n1766);
and gate_1748(n1768,n1725,n1767);
not gate_1749(n1769,n1768);
and gate_1750(n1770,n27,n1769);
not gate_1751(n1771,n1770);
and gate_1752(n1772,n25,n1695);
not gate_1753(n1773,n1772);
and gate_1754(n1774,pi4,n1737);
not gate_1755(n1775,n1774);
and gate_1756(n1776,n1773,n1775);
not gate_1757(n1777,n1776);
and gate_1758(n1778,n1022,n1777);
and gate_1759(n1779,n23,n1778);
not gate_1760(n1780,n1779);
and gate_1761(n1781,pi5,n1737);
not gate_1762(n1782,n1781);
and gate_1763(n1783,n1773,n1782);
not gate_1764(n1784,n1783);
and gate_1765(n1785,n24,n1784);
not gate_1766(n1786,n1785);
and gate_1767(n1787,n1021,n1674);
not gate_1768(n1788,n1787);
and gate_1769(n1789,n1786,n1788);
not gate_1770(n1790,n1789);
and gate_1771(n1791,pi3,n1790);
not gate_1772(n1792,n1791);
and gate_1773(n1793,n1780,n1792);
not gate_1774(n1794,n1793);
and gate_1775(n1795,pi9,n1794);
not gate_1776(n1796,n1795);
and gate_1777(n1797,n28,n100);
not gate_1778(n1798,n1797);
and gate_1779(n1799,n91,n1024);
not gate_1780(n1800,n1799);
and gate_1781(n1801,n1798,n1800);
and gate_1782(n1802,n173,n1801);
not gate_1783(n1803,n1802);
and gate_1784(n1804,n1796,n1803);
not gate_1785(n1805,n1804);
and gate_1786(n1806,pi2,n1805);
not gate_1787(n1807,n1806);
and gate_1788(n1808,n1687,n1691);
not gate_1789(n1809,n1808);
and gate_1790(n1810,n384,n1023);
and gate_1791(n1811,n1809,n1810);
and gate_1792(n1812,n23,n1811);
not gate_1793(n1813,n1812);
and gate_1794(n1814,n477,n995);
not gate_1795(n1815,n1814);
and gate_1796(n1816,n1813,n1815);
not gate_1797(n1817,n1816);
and gate_1798(n1818,pi6,n1817);
not gate_1799(n1819,n1818);
and gate_1800(n1820,pi3,n26);
not gate_1801(n1821,n1820);
and gate_1802(n1822,n384,n1808);
and gate_1803(n1823,n1020,n1822);
and gate_1804(n1824,n1820,n1823);
not gate_1805(n1825,n1824);
and gate_1806(n1826,n1819,n1825);
not gate_1807(n1827,n1826);
and gate_1808(n1828,n22,n1827);
not gate_1809(n1829,n1828);
and gate_1810(n1830,n1807,n1829);
not gate_1811(n1831,n1830);
and gate_1812(n1832,n21,n1831);
not gate_1813(n1833,n1832);
and gate_1814(n1834,n23,n99);
not gate_1815(n1835,n1834);
and gate_1816(n1836,pi3,n1625);
not gate_1817(n1837,n1836);
and gate_1818(n1838,n1835,n1837);
not gate_1819(n1839,n1838);
and gate_1820(n1840,pi2,n1839);
not gate_1821(n1841,n1840);
and gate_1822(n1842,n131,n1509);
not gate_1823(n1843,n1842);
and gate_1824(n1844,n1841,n1843);
not gate_1825(n1845,n1844);
and gate_1826(n1846,n29,n1845);
not gate_1827(n1847,n1846);
and gate_1828(n1848,pi3,n123);
not gate_1829(n1849,n1848);
and gate_1830(n1850,n22,n1848);
not gate_1831(n1851,n1850);
and gate_1832(n1852,n1847,n1851);
not gate_1833(n1853,n1852);
and gate_1834(n1854,pi4,n1853);
not gate_1835(n1855,n1854);
and gate_1836(n1856,n26,n952);
and gate_1837(n1857,pi2,n1856);
not gate_1838(n1858,n1857);
and gate_1839(n1859,n123,n131);
not gate_1840(n1860,n1859);
and gate_1841(n1861,n1858,n1860);
not gate_1842(n1862,n1861);
and gate_1843(n1863,n23,n1862);
not gate_1844(n1864,n1863);
and gate_1845(n1865,n288,n1279);
not gate_1846(n1866,n1865);
and gate_1847(n1867,n1864,n1866);
not gate_1848(n1868,n1867);
and gate_1849(n1869,n24,n1868);
not gate_1850(n1870,n1869);
and gate_1851(n1871,n1855,n1870);
not gate_1852(n1872,n1871);
and gate_1853(n1873,n28,n1872);
not gate_1854(n1874,n1873);
and gate_1855(n1875,pi5,n123);
not gate_1856(n1876,n1875);
and gate_1857(n1877,n1665,n1875);
not gate_1858(n1878,n1877);
and gate_1859(n1879,n23,n1625);
not gate_1860(n1880,n1879);
and gate_1861(n1881,n264,n1157);
not gate_1862(n1882,n1881);
and gate_1863(n1883,n1880,n1882);
not gate_1864(n1884,n1883);
and gate_1865(n1885,n1174,n1884);
not gate_1866(n1886,n1885);
and gate_1867(n1887,n1878,n1886);
not gate_1868(n1888,n1887);
and gate_1869(n1889,pi8,n1888);
not gate_1870(n1890,n1889);
and gate_1871(n1891,n1874,n1890);
not gate_1872(n1892,n1891);
and gate_1873(n1893,pi1,n1892);
not gate_1874(n1894,n1893);
and gate_1875(n1895,n1833,n1894);
not gate_1876(n1896,n1895);
and gate_1877(n1897,pi7,n1896);
not gate_1878(n1898,n1897);
and gate_1879(n1899,n1771,n1898);
not gate_1880(n1900,n1899);
and gate_1881(n1901,n20,n1900);
not gate_1882(n1902,n1901);
and gate_1883(n1903,n1664,n1902);
not gate_1884(po2,n1903);
and gate_1885(n1905,n20,n1476);
and gate_1886(n1906,n24,n949);
and gate_1887(n1907,n1905,n1906);
not gate_1888(n1908,n1907);
and gate_1889(n1909,pi0,n23);
not gate_1890(n1910,n1909);
and gate_1891(n1911,n587,n910);
not gate_1892(n1912,n1911);
and gate_1893(n1913,n979,n1912);
and gate_1894(n1914,n1909,n1913);
not gate_1895(n1915,n1914);
and gate_1896(n1916,n1908,n1915);
not gate_1897(n1917,n1916);
and gate_1898(n1918,n22,n1917);
not gate_1899(n1919,n1918);
and gate_1900(n1920,n785,n949);
and gate_1901(n1921,n1070,n1920);
not gate_1902(n1922,n1921);
and gate_1903(n1923,n1919,n1922);
not gate_1904(n1924,n1923);
and gate_1905(n1925,n26,n372);
not gate_1906(n1926,n1925);
and gate_1907(n1927,pi6,n232);
not gate_1908(n1928,n1927);
and gate_1909(n1929,n1926,n1928);
not gate_1910(n1930,n1929);
and gate_1911(n1931,n1924,n1930);
not gate_1912(n1932,n1931);
and gate_1913(n1933,n20,n131);
and gate_1914(n1934,n39,n1320);
and gate_1915(n1935,n1933,n1934);
not gate_1916(n1936,n1935);
and gate_1917(n1937,n26,n232);
and gate_1918(n1938,n889,n1937);
not gate_1919(n1939,n1938);
and gate_1920(n1940,n917,n1320);
not gate_1921(n1941,n1940);
and gate_1922(n1942,n1939,n1941);
not gate_1923(n1943,n1942);
and gate_1924(n1944,n535,n1943);
not gate_1925(n1945,n1944);
and gate_1926(n1946,n1936,n1945);
not gate_1927(n1947,n1946);
and gate_1928(n1948,pi1,n1947);
not gate_1929(n1949,n1948);
and gate_1930(n1950,n84,n917);
and gate_1931(n1951,n247,n1324);
and gate_1932(n1952,n1950,n1951);
not gate_1933(n1953,n1952);
and gate_1934(n1954,n1949,n1953);
not gate_1935(n1955,n1954);
and gate_1936(n1956,n1072,n1955);
not gate_1937(n1957,n1956);
and gate_1938(n1958,n1319,n1751);
not gate_1939(n1959,n1958);
and gate_1940(n1960,n1668,n1959);
and gate_1941(n1961,pi1,n1960);
not gate_1942(n1962,n1961);
and gate_1943(n1963,n21,n983);
and gate_1944(n1964,pi6,n39);
not gate_1945(n1965,n1964);
and gate_1946(n1966,n1963,n1964);
not gate_1947(n1967,n1966);
and gate_1948(n1968,n1962,n1967);
not gate_1949(n1969,n1968);
and gate_1950(n1970,n22,n1969);
not gate_1951(n1971,n1970);
and gate_1952(n1972,n39,n90);
and gate_1953(n1973,n1138,n1972);
not gate_1954(n1974,n1973);
and gate_1955(n1975,n1971,n1974);
not gate_1956(n1976,n1975);
and gate_1957(n1977,n20,n1976);
not gate_1958(n1978,n1977);
and gate_1959(n1979,n55,n74);
and gate_1960(n1980,n1972,n1979);
not gate_1961(n1981,n1980);
and gate_1962(n1982,n1978,n1981);
not gate_1963(n1983,n1982);
and gate_1964(n1984,n730,n1983);
not gate_1965(n1985,n1984);
and gate_1966(n1986,n927,n1197);
and gate_1967(n1987,n23,n1986);
not gate_1968(n1988,n1987);
and gate_1969(n1989,n25,n133);
not gate_1970(n1990,n1989);
and gate_1971(n1991,n1876,n1990);
not gate_1972(n1992,n1991);
and gate_1973(n1993,n1491,n1992);
not gate_1974(n1994,n1993);
and gate_1975(n1995,n1988,n1994);
not gate_1976(n1996,n1995);
and gate_1977(n1997,pi4,n1996);
not gate_1978(n1998,n1997);
and gate_1979(n1999,pi6,n188);
and gate_1980(n2000,pi3,n983);
and gate_1981(n2001,n1999,n2000);
not gate_1982(n2002,n2001);
and gate_1983(n2003,n1998,n2002);
not gate_1984(n2004,n2003);
and gate_1985(n2005,n21,n2004);
not gate_1986(n2006,n2005);
and gate_1987(n2007,n90,n190);
and gate_1988(n2008,n997,n2007);
not gate_1989(n2009,n2008);
and gate_1990(n2010,n2006,n2009);
not gate_1991(n2011,n2010);
and gate_1992(n2012,pi8,n2011);
not gate_1993(n2013,n2012);
and gate_1994(n2014,n1019,n1586);
not gate_1995(n2015,n2014);
and gate_1996(n2016,n26,n181);
and gate_1997(n2017,n1021,n2016);
not gate_1998(n2018,n2017);
and gate_1999(n2019,n2015,n2018);
not gate_2000(n2020,n2019);
and gate_2001(n2021,n354,n2020);
and gate_2002(n2022,pi1,n2021);
not gate_2003(n2023,n2022);
and gate_2004(n2024,n2013,n2023);
not gate_2005(n2025,n2024);
and gate_2006(n2026,pi0,n2025);
not gate_2007(n2027,n2026);
and gate_2008(n2028,n47,n1665);
and gate_2009(n2029,n69,n311);
and gate_2010(n2030,n2028,n2029);
not gate_2011(n2031,n2030);
and gate_2012(n2032,n2027,n2031);
and gate_2013(n2033,n424,n563);
and gate_2014(n2034,n1335,n2033);
not gate_2015(n2035,n2034);
and gate_2016(n2036,n564,n1299);
and gate_2017(n2037,n1668,n2036);
not gate_2018(n2038,n2037);
and gate_2019(n2039,n2035,n2038);
not gate_2020(n2040,n2039);
and gate_2021(n2041,pi3,n2040);
not gate_2022(n2042,n2041);
and gate_2023(n2043,n545,n1928);
not gate_2024(n2044,n2043);
and gate_2025(n2045,n1420,n2044);
and gate_2026(n2046,pi0,n2045);
not gate_2027(n2047,n2046);
and gate_2028(n2048,n47,n1937);
not gate_2029(n2049,n2048);
and gate_2030(n2050,n2047,n2049);
not gate_2031(n2051,n2050);
and gate_2032(n2052,n23,n2051);
not gate_2033(n2053,n2052);
and gate_2034(n2054,n2042,n2053);
not gate_2035(n2055,n2054);
and gate_2036(n2056,n25,n2055);
not gate_2037(n2057,n2056);
and gate_2038(n2058,n76,n1695);
not gate_2039(n2059,n2058);
and gate_2040(n2060,pi0,n1332);
not gate_2041(n2061,n2060);
and gate_2042(n2062,n1215,n2061);
not gate_2043(n2063,n2062);
and gate_2044(n2064,n28,n2063);
not gate_2045(n2065,n2064);
and gate_2046(n2066,n2059,n2065);
not gate_2047(n2067,n2066);
and gate_2048(n2068,n255,n2067);
not gate_2049(n2069,n2068);
and gate_2050(n2070,pi3,n2048);
not gate_2051(n2071,n2070);
and gate_2052(n2072,n2069,n2071);
not gate_2053(n2073,n2072);
and gate_2054(n2074,pi5,n2073);
not gate_2055(n2075,n2074);
and gate_2056(n2076,n2057,n2075);
not gate_2057(n2077,n2076);
and gate_2058(n2078,n29,n2077);
not gate_2059(n2079,n2078);
and gate_2060(n2080,pi5,n421);
and gate_2061(n2081,pi1,n2080);
not gate_2062(n2082,n2081);
and gate_2063(n2083,n26,n419);
and gate_2064(n2084,n350,n2083);
not gate_2065(n2085,n2084);
and gate_2066(n2086,n2082,n2085);
not gate_2067(n2087,n2086);
and gate_2068(n2088,n532,n1910);
not gate_2069(n2089,n2088);
and gate_2070(n2090,n2087,n2089);
not gate_2071(n2091,n2090);
and gate_2072(n2092,n25,pi8);
not gate_2073(n2093,n2092);
and gate_2074(n2094,n212,n2093);
not gate_2075(n2095,n2094);
and gate_2076(n2096,n20,pi8);
not gate_2077(n2097,n2096);
and gate_2078(n2098,pi0,n28);
not gate_2079(n2099,n2098);
and gate_2080(n2100,n2097,n2099);
not gate_2081(n2101,n2100);
and gate_2082(n2102,n2094,n2101);
and gate_2083(n2103,n1504,n2102);
not gate_2084(n2104,n2103);
and gate_2085(n2105,n1880,n2104);
not gate_2086(n2106,n2105);
and gate_2087(n2107,n27,n2106);
not gate_2088(n2108,n2107);
and gate_2089(n2109,n20,pi5);
not gate_2090(n2110,n2109);
and gate_2091(n2111,n1737,n2109);
not gate_2092(n2112,n2111);
and gate_2093(n2113,pi8,n1627);
and gate_2094(n2114,n2110,n2113);
not gate_2095(n2115,n2114);
and gate_2096(n2116,n2112,n2115);
not gate_2097(n2117,n2116);
and gate_2098(n2118,n255,n2117);
not gate_2099(n2119,n2118);
and gate_2100(n2120,n2108,n2119);
not gate_2101(n2121,n2120);
and gate_2102(n2122,n21,n2121);
not gate_2103(n2123,n2122);
and gate_2104(n2124,n25,n1740);
and gate_2105(n2125,pi0,n2124);
not gate_2106(n2126,n2125);
and gate_2107(n2127,n1668,n2109);
not gate_2108(n2128,n2127);
and gate_2109(n2129,n2126,n2128);
not gate_2110(n2130,n2129);
and gate_2111(n2131,pi1,n255);
not gate_2112(n2132,n2131);
and gate_2113(n2133,n2130,n2131);
not gate_2114(n2134,n2133);
and gate_2115(n2135,n2123,n2134);
and gate_2116(n2136,n2091,n2135);
not gate_2117(n2137,n2136);
and gate_2118(n2138,pi9,n2137);
not gate_2119(n2139,n2138);
and gate_2120(n2140,n2079,n2139);
not gate_2121(n2141,n2140);
and gate_2122(n2142,pi2,n2141);
not gate_2123(n2143,n2142);
and gate_2124(n2144,n42,n478);
not gate_2125(n2145,n2144);
and gate_2126(n2146,n70,n2145);
and gate_2127(n2147,n20,n2146);
not gate_2128(n2148,n2147);
and gate_2129(n2149,n32,n69);
not gate_2130(n2150,n2149);
and gate_2131(n2151,n196,n1127);
not gate_2132(n2152,n2151);
and gate_2133(n2153,n2150,n2152);
not gate_2134(n2154,n2153);
and gate_2135(n2155,pi0,n2154);
not gate_2136(n2156,n2155);
and gate_2137(n2157,n2148,n2156);
not gate_2138(n2158,n2157);
and gate_2139(n2159,n27,n2158);
not gate_2140(n2160,n2159);
and gate_2141(n2161,n20,n25);
not gate_2142(n2162,n2161);
and gate_2143(n2163,n164,n2162);
not gate_2144(n2164,n2163);
and gate_2145(n2165,n204,n2163);
and gate_2146(n2166,n195,n2165);
and gate_2147(n2167,n1197,n2166);
not gate_2148(n2168,n2167);
and gate_2149(n2169,n2160,n2168);
not gate_2150(n2170,n2169);
and gate_2151(n2171,pi3,n2170);
not gate_2152(n2172,n2171);
and gate_2153(n2173,n69,n232);
not gate_2154(n2174,n2173);
and gate_2155(n2175,n90,n424);
not gate_2156(n2176,n2175);
and gate_2157(n2177,n2174,n2176);
not gate_2158(n2178,n2177);
and gate_2159(n2179,n20,n2178);
not gate_2160(n2180,n2179);
and gate_2161(n2181,pi0,n25);
and gate_2162(n2182,pi6,n372);
and gate_2163(n2183,n2181,n2182);
not gate_2164(n2184,n2183);
and gate_2165(n2185,n2180,n2184);
not gate_2166(n2186,n2185);
and gate_2167(n2187,pi9,n2186);
not gate_2168(n2188,n2187);
and gate_2169(n2189,n20,n1625);
and gate_2170(n2190,n311,n2189);
not gate_2171(n2191,n2190);
and gate_2172(n2192,n2188,n2191);
not gate_2173(n2193,n2192);
and gate_2174(n2194,n23,n2193);
not gate_2175(n2195,n2194);
and gate_2176(n2196,n2172,n2195);
not gate_2177(n2197,n2196);
and gate_2178(n2198,pi1,n2197);
not gate_2179(n2199,n2198);
and gate_2180(n2200,pi3,n1402);
not gate_2181(n2201,n2200);
and gate_2182(n2202,n190,n1506);
not gate_2183(n2203,n2202);
and gate_2184(n2204,n2201,n2203);
not gate_2185(n2205,n2204);
and gate_2186(n2206,pi5,n2205);
not gate_2187(n2207,n2206);
and gate_2188(n2208,n124,n153);
and gate_2189(n2209,n23,n2208);
not gate_2190(n2210,n2209);
and gate_2191(n2211,n2207,n2210);
not gate_2192(n2212,n2211);
and gate_2193(n2213,pi0,n2212);
not gate_2194(n2214,n2213);
and gate_2195(n2215,n841,n1715);
not gate_2196(n2216,n2215);
and gate_2197(n2217,n181,n2216);
and gate_2198(n2218,n20,n2217);
not gate_2199(n2219,n2218);
and gate_2200(n2220,n2214,n2219);
not gate_2201(n2221,n2220);
and gate_2202(n2222,pi8,n2221);
not gate_2203(n2223,n2222);
and gate_2204(n2224,n26,n32);
not gate_2205(n2225,n2224);
and gate_2206(n2226,n1299,n2162);
and gate_2207(n2227,n2224,n2226);
and gate_2208(n2228,pi3,n2227);
not gate_2209(n2229,n2228);
and gate_2210(n2230,n2223,n2229);
not gate_2211(n2231,n2230);
and gate_2212(n2232,n21,n2231);
not gate_2213(n2233,n2232);
and gate_2214(n2234,n2199,n2233);
not gate_2215(n2235,n2234);
and gate_2216(n2236,n22,n2235);
not gate_2217(n2237,n2236);
and gate_2218(n2238,n2143,n2237);
not gate_2219(n2239,n2238);
and gate_2220(n2240,n24,n2239);
not gate_2221(n2241,n2240);
and gate_2222(n2242,n21,n32);
not gate_2223(n2243,n2242);
and gate_2224(n2244,pi1,n424);
not gate_2225(n2245,n2244);
and gate_2226(n2246,n21,n423);
not gate_2227(n2247,n2246);
and gate_2228(n2248,n2245,n2247);
and gate_2229(n2249,n29,n2248);
not gate_2230(n2250,n2249);
and gate_2231(n2251,n2243,n2250);
not gate_2232(n2252,n2251);
and gate_2233(n2253,pi5,n2252);
not gate_2234(n2254,n2253);
and gate_2235(n2255,n477,n1480);
not gate_2236(n2256,n2255);
and gate_2237(n2257,n2254,n2256);
not gate_2238(n2258,n2257);
and gate_2239(n2259,pi3,n2258);
not gate_2240(n2260,n2259);
and gate_2241(n2261,n204,n701);
not gate_2242(n2262,n2261);
and gate_2243(n2263,n50,n2262);
and gate_2244(n2264,n605,n2263);
not gate_2245(n2265,n2264);
and gate_2246(n2266,n2260,n2265);
not gate_2247(n2267,n2266);
and gate_2248(n2268,n22,n2267);
not gate_2249(n2269,n2268);
and gate_2250(n2270,n21,n1491);
not gate_2251(n2271,n2270);
and gate_2252(n2272,n2132,n2271);
not gate_2253(n2273,n2272);
and gate_2254(n2274,n462,n2273);
not gate_2255(n2275,n2274);
and gate_2256(n2276,pi7,n39);
and gate_2257(n2277,n1476,n2276);
not gate_2258(n2278,n2277);
and gate_2259(n2279,n2275,n2278);
not gate_2260(n2280,n2279);
and gate_2261(n2281,n25,n2280);
not gate_2262(n2282,n2281);
and gate_2263(n2283,pi1,n436);
not gate_2264(n2284,n2283);
and gate_2265(n2285,n2282,n2284);
not gate_2266(n2286,n2285);
and gate_2267(n2287,pi2,n2286);
not gate_2268(n2288,n2287);
and gate_2269(n2289,n2269,n2288);
not gate_2270(n2290,n2289);
and gate_2271(n2291,n20,n2290);
not gate_2272(n2292,n2291);
and gate_2273(n2293,n192,n858);
and gate_2274(n2294,n1912,n2293);
and gate_2275(n2295,pi2,n2294);
not gate_2276(n2296,n2295);
and gate_2277(n2297,pi3,n181);
not gate_2278(n2298,n2297);
and gate_2279(n2299,n407,n2298);
not gate_2280(n2300,n2299);
and gate_2281(n2301,n337,n2300);
not gate_2282(n2302,n2301);
and gate_2283(n2303,n2296,n2302);
not gate_2284(n2304,n2303);
and gate_2285(n2305,n25,n2304);
not gate_2286(n2306,n2305);
and gate_2287(n2307,n22,n121);
and gate_2288(n2308,n1477,n2272);
not gate_2289(n2309,n2308);
and gate_2290(n2310,n2307,n2309);
not gate_2291(n2311,n2310);
and gate_2292(n2312,n2306,n2311);
not gate_2293(n2313,n2312);
and gate_2294(n2314,n28,n2313);
not gate_2295(n2315,n2314);
and gate_2296(n2316,n305,n1114);
not gate_2297(n2317,n2316);
and gate_2298(n2318,n265,n338);
not gate_2299(n2319,n2318);
and gate_2300(n2320,n2317,n2319);
and gate_2301(n2321,n27,n2320);
not gate_2302(n2322,n2321);
and gate_2303(n2323,pi1,n727);
and gate_2304(n2324,n466,n2323);
not gate_2305(n2325,n2324);
and gate_2306(n2326,n2322,n2325);
not gate_2307(n2327,n2326);
and gate_2308(n2328,pi9,n2327);
not gate_2309(n2329,n2328);
and gate_2310(n2330,pi2,n190);
not gate_2311(n2331,n2330);
and gate_2312(n2332,n264,n2330);
not gate_2313(n2333,n2332);
and gate_2314(n2334,n2329,n2333);
not gate_2315(n2335,n2334);
and gate_2316(n2336,pi8,n2335);
not gate_2317(n2337,n2336);
and gate_2318(n2338,n2315,n2337);
not gate_2319(n2339,n2338);
and gate_2320(n2340,pi0,n2339);
not gate_2321(n2341,n2340);
and gate_2322(n2342,n2292,n2341);
not gate_2323(n2343,n2342);
and gate_2324(n2344,n26,n2343);
not gate_2325(n2345,n2344);
and gate_2326(n2346,n563,n1299);
and gate_2327(n2347,n426,n2346);
and gate_2328(n2348,n22,n2347);
not gate_2329(n2349,n2348);
and gate_2330(n2350,pi7,n2163);
not gate_2331(n2351,n2350);
and gate_2332(n2352,n351,n545);
not gate_2333(n2353,n2352);
and gate_2334(n2354,n2351,n2353);
and gate_2335(n2355,pi2,n2354);
not gate_2336(n2356,n2355);
and gate_2337(n2357,n2349,n2356);
not gate_2338(n2358,n2357);
and gate_2339(n2359,pi3,n2358);
not gate_2340(n2360,n2359);
and gate_2341(n2361,n37,n154);
and gate_2342(n2362,n76,n2361);
not gate_2343(n2363,n2362);
and gate_2344(n2364,n2360,n2363);
not gate_2345(n2365,n2364);
and gate_2346(n2366,n28,n2365);
not gate_2347(n2367,n2366);
and gate_2348(n2368,n47,n840);
not gate_2349(n2369,n2368);
and gate_2350(n2370,n351,n371);
not gate_2351(n2371,n2370);
and gate_2352(n2372,n1909,n2371);
not gate_2353(n2373,n2372);
and gate_2354(n2374,n2369,n2373);
not gate_2355(n2375,n2374);
and gate_2356(n2376,pi2,n2375);
not gate_2357(n2377,n2376);
and gate_2358(n2378,n22,n264);
not gate_2359(n2379,n2378);
and gate_2360(n2380,n76,n2378);
not gate_2361(n2381,n2380);
and gate_2362(n2382,n2377,n2381);
not gate_2363(n2383,n2382);
and gate_2364(n2384,n372,n2383);
not gate_2365(n2385,n2384);
and gate_2366(n2386,n2367,n2385);
not gate_2367(n2387,n2386);
and gate_2368(n2388,pi9,n2387);
not gate_2369(n2389,n2388);
and gate_2370(n2390,n20,n772);
not gate_2371(n2391,n2390);
and gate_2372(n2392,pi0,n633);
not gate_2373(n2393,n2392);
and gate_2374(n2394,n424,n2392);
not gate_2375(n2395,n2394);
and gate_2376(n2396,n2391,n2395);
not gate_2377(n2397,n2396);
and gate_2378(n2398,n23,n2397);
not gate_2379(n2399,n2398);
and gate_2380(n2400,n22,n421);
not gate_2381(n2401,n2400);
and gate_2382(n2402,n531,n2400);
not gate_2383(n2403,n2402);
and gate_2384(n2404,n2399,n2403);
not gate_2385(n2405,n2404);
and gate_2386(n2406,n25,n2405);
not gate_2387(n2407,n2406);
and gate_2388(n2408,pi5,n232);
and gate_2389(n2409,n20,n30);
and gate_2390(n2410,n2408,n2409);
not gate_2391(n2411,n2410);
and gate_2392(n2412,n2407,n2411);
not gate_2393(n2413,n2412);
and gate_2394(n2414,n580,n2413);
not gate_2395(n2415,n2414);
and gate_2396(n2416,n2389,n2415);
not gate_2397(n2417,n2416);
and gate_2398(n2418,pi6,n2417);
not gate_2399(n2419,n2418);
and gate_2400(n2420,n2345,n2419);
not gate_2401(n2421,n2420);
and gate_2402(n2422,pi4,n2421);
not gate_2403(n2423,n2422);
and gate_2404(n2424,n2241,n2423);
and gate_2405(n2425,n2032,n2424);
and gate_2406(n2426,n1985,n2425);
and gate_2407(n2427,n1957,n2426);
and gate_2408(n2428,n1932,n2427);
not gate_2409(po3,n2428);
and gate_2410(n2430,pi3,pi4);
not gate_2411(n2431,n2430);
and gate_2412(n2432,n1666,n2431);
not gate_2413(n2433,n2432);
and gate_2414(n2434,n364,n2432);
and gate_2415(n2435,n730,n2434);
and gate_2416(n2436,n1695,n2435);
and gate_2417(n2437,pi0,n2436);
not gate_2418(n2438,n2437);
and gate_2419(n2439,n20,n37);
and gate_2420(n2440,n419,n1152);
and gate_2421(n2441,n2439,n2440);
not gate_2422(n2442,n2441);
and gate_2423(n2443,n2438,n2442);
not gate_2424(n2444,n2443);
and gate_2425(n2445,n927,n2444);
not gate_2426(n2446,n2445);
and gate_2427(n2447,n239,n662);
not gate_2428(n2448,n2447);
and gate_2429(n2449,pi0,n858);
not gate_2430(n2450,n2449);
and gate_2431(n2451,n925,n2449);
not gate_2432(n2452,n2451);
and gate_2433(n2453,n2448,n2452);
not gate_2434(n2454,n2453);
and gate_2435(n2455,n27,n2454);
not gate_2436(n2456,n2455);
and gate_2437(n2457,n408,n690);
not gate_2438(n2458,n2457);
and gate_2439(n2459,n2456,n2458);
not gate_2440(n2460,n2459);
and gate_2441(n2461,n24,n2460);
not gate_2442(n2462,n2461);
and gate_2443(n2463,pi0,n37);
and gate_2444(n2464,pi4,n190);
and gate_2445(n2465,n2463,n2464);
not gate_2446(n2466,n2465);
and gate_2447(n2467,n2462,n2466);
not gate_2448(n2468,n2467);
and gate_2449(n2469,pi8,n2468);
not gate_2450(n2470,n2469);
and gate_2451(n2471,n20,n874);
and gate_2452(n2472,n32,n1421);
and gate_2453(n2473,n2471,n2472);
not gate_2454(n2474,n2473);
and gate_2455(n2475,n2470,n2474);
not gate_2456(n2476,n2475);
and gate_2457(n2477,n1628,n2476);
not gate_2458(n2478,n2477);
and gate_2459(n2479,pi3,n196);
not gate_2460(n2480,n2479);
and gate_2461(n2481,n32,n842);
not gate_2462(n2482,n2481);
and gate_2463(n2483,n2480,n2482);
not gate_2464(n2484,n2483);
and gate_2465(n2485,n26,n2484);
not gate_2466(n2486,n2485);
and gate_2467(n2487,n1128,n2094);
and gate_2468(n2488,n357,n2487);
not gate_2469(n2489,n2488);
and gate_2470(n2490,n2486,n2489);
not gate_2471(n2491,n2490);
and gate_2472(n2492,n27,n2491);
not gate_2473(n2493,n2492);
and gate_2474(n2494,n124,n134);
not gate_2475(n2495,n2494);
and gate_2476(n2496,n962,n2494);
and gate_2477(n2497,n950,n2496);
and gate_2478(n2498,pi8,n2497);
not gate_2479(n2499,n2498);
and gate_2480(n2500,n25,n1737);
and gate_2481(n2501,n23,n2500);
not gate_2482(n2502,n2501);
and gate_2483(n2503,n2499,n2502);
not gate_2484(n2504,n2503);
and gate_2485(n2505,pi7,n2504);
not gate_2486(n2506,n2505);
and gate_2487(n2507,n2493,n2506);
not gate_2488(n2508,n2507);
and gate_2489(n2509,n24,n2508);
not gate_2490(n2510,n2509);
and gate_2491(n2511,n305,n355);
and gate_2492(n2512,n279,n2511);
and gate_2493(n2513,n26,n2512);
not gate_2494(n2514,n2513);
and gate_2495(n2515,pi6,n278);
and gate_2496(n2516,n304,n2515);
not gate_2497(n2517,n2516);
and gate_2498(n2518,n2514,n2517);
not gate_2499(n2519,n2518);
and gate_2500(n2520,n27,n2519);
not gate_2501(n2521,n2520);
and gate_2502(n2522,n357,n1293);
and gate_2503(n2523,n25,n2522);
not gate_2504(n2524,n2523);
and gate_2505(n2525,n2521,n2524);
not gate_2506(n2526,n2525);
and gate_2507(n2527,pi4,n2526);
not gate_2508(n2528,n2527);
and gate_2509(n2529,n2510,n2528);
not gate_2510(n2530,n2529);
and gate_2511(n2531,pi2,n2530);
not gate_2512(n2532,n2531);
and gate_2513(n2533,n26,n188);
not gate_2514(n2534,n2533);
and gate_2515(n2535,n322,n2534);
not gate_2516(n2536,n2535);
and gate_2517(n2537,n70,n2536);
and gate_2518(n2538,pi4,n2537);
not gate_2519(n2539,n2538);
and gate_2520(n2540,n1601,n2539);
not gate_2521(n2541,n2540);
and gate_2522(n2542,n28,n2541);
not gate_2523(n2543,n2542);
and gate_2524(n2544,n189,n2494);
and gate_2525(n2545,n122,n2544);
and gate_2526(n2546,n1686,n2545);
not gate_2527(n2547,n2546);
and gate_2528(n2548,n2543,n2547);
not gate_2529(n2549,n2548);
and gate_2530(n2550,n23,n2549);
not gate_2531(n2551,n2550);
and gate_2532(n2552,n24,n27);
not gate_2533(n2553,n2552);
and gate_2534(n2554,n140,n2553);
and gate_2535(n2555,n2093,n2554);
not gate_2536(n2556,n2555);
and gate_2537(n2557,n212,n1422);
not gate_2538(n2558,n2557);
and gate_2539(n2559,n2556,n2558);
and gate_2540(n2560,pi6,n2559);
not gate_2541(n2561,n2560);
and gate_2542(n2562,n1021,n1925);
not gate_2543(n2563,n2562);
and gate_2544(n2564,n2561,n2563);
not gate_2545(n2565,n2564);
and gate_2546(n2566,n29,n2565);
not gate_2547(n2567,n2566);
and gate_2548(n2568,n32,n1453);
and gate_2549(n2569,n1019,n2568);
not gate_2550(n2570,n2569);
and gate_2551(n2571,n2567,n2570);
not gate_2552(n2572,n2571);
and gate_2553(n2573,pi3,n2572);
not gate_2554(n2574,n2573);
and gate_2555(n2575,n2551,n2574);
not gate_2556(n2576,n2575);
and gate_2557(n2577,n22,n2576);
not gate_2558(n2578,n2577);
and gate_2559(n2579,n2532,n2578);
not gate_2560(n2580,n2579);
and gate_2561(n2581,pi0,n2580);
not gate_2562(n2582,n2581);
and gate_2563(n2583,pi2,n149);
not gate_2564(n2584,n2583);
and gate_2565(n2585,n154,n2584);
not gate_2566(n2586,n2585);
and gate_2567(n2587,n28,n2586);
not gate_2568(n2588,n2587);
and gate_2569(n2589,n2401,n2588);
not gate_2570(n2590,n2589);
and gate_2571(n2591,pi4,n2590);
not gate_2572(n2592,n2591);
and gate_2573(n2593,n27,n2095);
and gate_2574(n2594,n165,n2593);
not gate_2575(n2595,n2594);
and gate_2576(n2596,n2592,n2595);
not gate_2577(n2597,n2596);
and gate_2578(n2598,pi6,n2597);
not gate_2579(n2599,n2598);
and gate_2580(n2600,n156,n2584);
not gate_2581(n2601,n2600);
and gate_2582(n2602,n1695,n2601);
not gate_2583(n2603,n2602);
and gate_2584(n2604,n2599,n2603);
not gate_2585(n2605,n2604);
and gate_2586(n2606,n29,n2605);
not gate_2587(n2607,n2606);
and gate_2588(n2608,pi4,n1937);
not gate_2589(n2609,n2608);
and gate_2590(n2610,n1019,n2182);
not gate_2591(n2611,n2610);
and gate_2592(n2612,n2609,n2611);
not gate_2593(n2613,n2612);
and gate_2594(n2614,pi2,n2613);
not gate_2595(n2615,n2614);
and gate_2596(n2616,n22,n1019);
and gate_2597(n2617,n26,n421);
not gate_2598(n2618,n2617);
and gate_2599(n2619,n2616,n2617);
not gate_2600(n2620,n2619);
and gate_2601(n2621,n2615,n2620);
not gate_2602(n2622,n2621);
and gate_2603(n2623,pi9,n2622);
not gate_2604(n2624,n2623);
and gate_2605(n2625,n2607,n2624);
not gate_2606(n2626,n2625);
and gate_2607(n2627,pi3,n2626);
not gate_2608(n2628,n2627);
and gate_2609(n2629,n69,n700);
not gate_2610(n2630,n2629);
and gate_2611(n2631,pi6,n426);
and gate_2612(n2632,n194,n312);
not gate_2613(n2633,n2632);
and gate_2614(n2634,n2631,n2633);
not gate_2615(n2635,n2634);
and gate_2616(n2636,n2630,n2635);
not gate_2617(n2637,n2636);
and gate_2618(n2638,pi4,n2637);
not gate_2619(n2639,n2638);
and gate_2620(n2640,n49,n278);
not gate_2621(n2641,n2640);
and gate_2622(n2642,n191,n320);
not gate_2623(n2643,n2642);
and gate_2624(n2644,n28,n2643);
not gate_2625(n2645,n2644);
and gate_2626(n2646,n2641,n2645);
not gate_2627(n2647,n2646);
and gate_2628(n2648,n26,n2647);
not gate_2629(n2649,n2648);
and gate_2630(n2650,pi7,n32);
and gate_2631(n2651,n99,n2650);
not gate_2632(n2652,n2651);
and gate_2633(n2653,n2649,n2652);
not gate_2634(n2654,n2653);
and gate_2635(n2655,n24,n2654);
not gate_2636(n2656,n2655);
and gate_2637(n2657,n2639,n2656);
not gate_2638(n2658,n2657);
and gate_2639(n2659,n874,n2658);
not gate_2640(n2660,n2659);
and gate_2641(n2661,n2628,n2660);
not gate_2642(n2662,n2661);
and gate_2643(n2663,n20,n2662);
not gate_2644(n2664,n2663);
and gate_2645(n2665,n2582,n2664);
and gate_2646(n2666,n2478,n2665);
and gate_2647(n2667,n2446,n2666);
not gate_2648(n2668,n2667);
and gate_2649(n2669,pi1,n2668);
not gate_2650(n2670,n2669);
and gate_2651(n2671,n926,n2094);
and gate_2652(n2672,n1628,n2671);
and gate_2653(n2673,pi3,n2672);
not gate_2654(n2674,n2673);
and gate_2655(n2675,n842,n1123);
not gate_2656(n2676,n2675);
and gate_2657(n2677,n2674,n2676);
not gate_2658(n2678,n2677);
and gate_2659(n2679,pi0,n2678);
not gate_2660(n2680,n2679);
and gate_2661(n2681,n20,n304);
and gate_2662(n2682,n34,n2681);
not gate_2663(n2683,n2682);
and gate_2664(n2684,n2680,n2683);
not gate_2665(n2685,n2684);
and gate_2666(n2686,n27,n2685);
not gate_2667(n2687,n2686);
and gate_2668(n2688,n1821,n1835);
not gate_2669(n2689,n2688);
and gate_2670(n2690,n20,n2276);
not gate_2671(n2691,n2690);
and gate_2672(n2692,n2689,n2690);
not gate_2673(n2693,n2692);
and gate_2674(n2694,n2687,n2693);
not gate_2675(n2695,n2694);
and gate_2676(n2696,n83,n2695);
not gate_2677(n2697,n2696);
and gate_2678(n2698,n166,n1691);
and gate_2679(n2699,pi0,n2698);
not gate_2680(n2700,n2699);
and gate_2681(n2701,pi7,n1235);
and gate_2682(n2702,n1809,n2701);
not gate_2683(n2703,n2702);
and gate_2684(n2704,n2700,n2703);
not gate_2685(n2705,n2704);
and gate_2686(n2706,n25,n2705);
not gate_2687(n2707,n2706);
and gate_2688(n2708,n24,n1197);
not gate_2689(n2709,n2708);
and gate_2690(n2710,n1422,n2709);
not gate_2691(n2711,n2710);
and gate_2692(n2712,n205,n2711);
and gate_2693(n2713,pi0,n2712);
not gate_2694(n2714,n2713);
and gate_2695(n2715,n2707,n2714);
not gate_2696(n2716,n2715);
and gate_2697(n2717,n23,n2716);
not gate_2698(n2718,n2717);
and gate_2699(n2719,pi0,n1809);
not gate_2700(n2720,n2719);
and gate_2701(n2721,n20,n1706);
not gate_2702(n2722,n2721);
and gate_2703(n2723,n2720,n2722);
not gate_2704(n2724,n2723);
and gate_2705(n2725,pi5,n2724);
not gate_2706(n2726,n2725);
and gate_2707(n2727,n1292,n2092);
not gate_2708(n2728,n2727);
and gate_2709(n2729,n2726,n2728);
not gate_2710(n2730,n2729);
and gate_2711(n2731,n26,n2730);
not gate_2712(n2732,n2731);
and gate_2713(n2733,n20,n24);
not gate_2714(n2734,n2733);
and gate_2715(n2735,n2500,n2733);
not gate_2716(n2736,n2735);
and gate_2717(n2737,n2732,n2736);
not gate_2718(n2738,n2737);
and gate_2719(n2739,n27,n2738);
not gate_2720(n2740,n2739);
and gate_2721(n2741,pi5,n1197);
and gate_2722(n2742,n2101,n2741);
and gate_2723(n2743,pi4,n2742);
not gate_2724(n2744,n2743);
and gate_2725(n2745,n2740,n2744);
not gate_2726(n2746,n2745);
and gate_2727(n2747,pi3,n2746);
not gate_2728(n2748,n2747);
and gate_2729(n2749,n2718,n2748);
not gate_2730(n2750,n2749);
and gate_2731(n2751,n22,n2750);
not gate_2732(n2752,n2751);
and gate_2733(n2753,pi0,n1509);
not gate_2734(n2754,n2753);
and gate_2735(n2755,n20,n1820);
not gate_2736(n2756,n2755);
and gate_2737(n2757,n2754,n2756);
not gate_2738(n2758,n2757);
and gate_2739(n2759,n24,n2758);
not gate_2740(n2760,n2759);
and gate_2741(n2761,n20,n23);
and gate_2742(n2762,n1152,n2761);
not gate_2743(n2763,n2762);
and gate_2744(n2764,n2760,n2763);
not gate_2745(n2765,n2764);
and gate_2746(n2766,n28,n2765);
not gate_2747(n2767,n2766);
and gate_2748(n2768,pi0,n1697);
not gate_2749(n2769,n2768);
and gate_2750(n2770,n2767,n2769);
not gate_2751(n2771,n2770);
and gate_2752(n2772,pi7,n2771);
not gate_2753(n2773,n2772);
and gate_2754(n2774,pi0,pi3);
not gate_2755(n2775,n2774);
and gate_2756(n2776,n166,n1707);
and gate_2757(n2777,n2774,n2776);
not gate_2758(n2778,n2777);
and gate_2759(n2779,n2773,n2778);
not gate_2760(n2780,n2779);
and gate_2761(n2781,pi5,n2780);
not gate_2762(n2782,n2781);
and gate_2763(n2783,n23,n1690);
not gate_2764(n2784,n2783);
and gate_2765(n2785,n1423,n1687);
and gate_2766(n2786,n2784,n2785);
and gate_2767(n2787,n20,n2786);
not gate_2768(n2788,n2787);
and gate_2769(n2789,pi4,n372);
and gate_2770(n2790,n1909,n2789);
not gate_2771(n2791,n2790);
and gate_2772(n2792,n2788,n2791);
not gate_2773(n2793,n2792);
and gate_2774(n2794,n69,n2793);
not gate_2775(n2795,n2794);
and gate_2776(n2796,n2782,n2795);
not gate_2777(n2797,n2796);
and gate_2778(n2798,pi2,n2797);
not gate_2779(n2799,n2798);
and gate_2780(n2800,n2752,n2799);
not gate_2781(n2801,n2800);
and gate_2782(n2802,pi9,n2801);
not gate_2783(n2803,n2802);
and gate_2784(n2804,n372,n1510);
not gate_2785(n2805,n2804);
and gate_2786(n2806,pi2,n1200);
and gate_2787(n2807,n1739,n2806);
not gate_2788(n2808,n2807);
and gate_2789(n2809,n2805,n2808);
not gate_2790(n2810,n2809);
and gate_2791(n2811,n24,n2810);
not gate_2792(n2812,n2811);
and gate_2793(n2813,n74,n1937);
not gate_2794(n2814,n2813);
and gate_2795(n2815,n2812,n2814);
not gate_2796(n2816,n2815);
and gate_2797(n2817,pi5,n2816);
not gate_2798(n2818,n2817);
and gate_2799(n2819,n421,n1154);
not gate_2800(n2820,n2819);
and gate_2801(n2821,n1320,n1687);
not gate_2802(n2822,n2821);
and gate_2803(n2823,n2820,n2822);
not gate_2804(n2824,n2823);
and gate_2805(n2825,n917,n2824);
not gate_2806(n2826,n2825);
and gate_2807(n2827,n2818,n2826);
not gate_2808(n2828,n2827);
and gate_2809(n2829,n20,n2828);
not gate_2810(n2830,n2829);
and gate_2811(n2831,pi6,n419);
not gate_2812(n2832,n2831);
and gate_2813(n2833,n2618,n2832);
not gate_2814(n2834,n2833);
and gate_2815(n2835,pi5,n2834);
and gate_2816(n2836,pi4,n2835);
not gate_2817(n2837,n2836);
and gate_2818(n2838,n983,n2182);
not gate_2819(n2839,n2838);
and gate_2820(n2840,n2837,n2839);
not gate_2821(n2841,n2840);
and gate_2822(n2842,pi2,n2841);
not gate_2823(n2843,n2842);
and gate_2824(n2844,n1616,n2831);
not gate_2825(n2845,n2844);
and gate_2826(n2846,n2843,n2845);
not gate_2827(n2847,n2846);
and gate_2828(n2848,pi0,n2847);
not gate_2829(n2849,n2848);
and gate_2830(n2850,n2830,n2849);
not gate_2831(n2851,n2850);
and gate_2832(n2852,pi3,n2851);
not gate_2833(n2853,n2852);
and gate_2834(n2854,n24,n1930);
not gate_2835(n2855,n2854);
and gate_2836(n2856,n372,n1152);
not gate_2837(n2857,n2856);
and gate_2838(n2858,n2855,n2857);
not gate_2839(n2859,n2858);
and gate_2840(n2860,n22,n2859);
not gate_2841(n2861,n2860);
and gate_2842(n2862,n82,n424);
and gate_2843(n2863,n1236,n2862);
not gate_2844(n2864,n2863);
and gate_2845(n2865,n2861,n2864);
not gate_2846(n2866,n2865);
and gate_2847(n2867,n25,n2866);
not gate_2848(n2868,n2867);
and gate_2849(n2869,n698,n1324);
not gate_2850(n2870,n2869);
and gate_2851(n2871,n24,n1452);
and gate_2852(n2872,n359,n2871);
not gate_2853(n2873,n2872);
and gate_2854(n2874,n2870,n2873);
not gate_2855(n2875,n2874);
and gate_2856(n2876,n211,n2875);
not gate_2857(n2877,n2876);
and gate_2858(n2878,n2868,n2877);
not gate_2859(n2879,n2878);
and gate_2860(n2880,n1909,n2879);
not gate_2861(n2881,n2880);
and gate_2862(n2882,n2853,n2881);
not gate_2863(n2883,n2882);
and gate_2864(n2884,n29,n2883);
not gate_2865(n2885,n2884);
and gate_2866(n2886,n2803,n2885);
and gate_2867(n2887,n2697,n2886);
not gate_2868(n2888,n2887);
and gate_2869(n2889,n21,n2888);
not gate_2870(n2890,n2889);
and gate_2871(n2891,n2670,n2890);
not gate_2872(po4,n2891);
and gate_2873(n2893,n232,n1154);
and gate_2874(n2894,n2471,n2893);
not gate_2875(n2895,n2894);
and gate_2876(n2896,n232,n874);
not gate_2877(n2897,n2896);
and gate_2878(n2898,n375,n2897);
not gate_2879(n2899,n2898);
and gate_2880(n2900,pi0,n2899);
not gate_2881(n2901,n2900);
and gate_2882(n2902,n592,n690);
not gate_2883(n2903,n2902);
and gate_2884(n2904,n2901,n2903);
not gate_2885(n2905,n2904);
and gate_2886(n2906,n1152,n2905);
not gate_2887(n2907,n2906);
and gate_2888(n2908,n2895,n2907);
not gate_2889(n2909,n2908);
and gate_2890(n2910,pi1,n2909);
not gate_2891(n2911,n2910);
and gate_2892(n2912,n84,n288);
and gate_2893(n2913,n106,n421);
and gate_2894(n2914,n2912,n2913);
not gate_2895(n2915,n2914);
and gate_2896(n2916,n2911,n2915);
not gate_2897(n2917,n2916);
and gate_2898(n2918,n952,n2917);
not gate_2899(n2919,n2918);
and gate_2900(n2920,pi6,n421);
and gate_2901(n2921,pi1,n983);
and gate_2902(n2922,n2920,n2921);
not gate_2903(n2923,n2922);
and gate_2904(n2924,n21,n979);
and gate_2905(n2925,n2083,n2924);
not gate_2906(n2926,n2925);
and gate_2907(n2927,n2923,n2926);
not gate_2908(n2928,n2927);
and gate_2909(n2929,n22,n2928);
and gate_2910(n2930,pi0,n2929);
not gate_2911(n2931,n2930);
and gate_2912(n2932,n76,n80);
and gate_2913(n2933,n372,n1625);
and gate_2914(n2934,n2932,n2933);
not gate_2915(n2935,n2934);
and gate_2916(n2936,n2931,n2935);
not gate_2917(n2937,n2936);
and gate_2918(n2938,n23,n2937);
not gate_2919(n2939,n2938);
and gate_2920(n2940,n712,n1695);
not gate_2921(n2941,n2940);
and gate_2922(n2942,n2391,n2941);
not gate_2923(n2943,n2942);
and gate_2924(n2944,n51,n2943);
and gate_2925(n2945,n522,n2944);
not gate_2926(n2946,n2945);
and gate_2927(n2947,n2939,n2946);
and gate_2928(n2948,n47,n504);
not gate_2929(n2949,n2948);
and gate_2930(n2950,n55,n506);
not gate_2931(n2951,n2950);
and gate_2932(n2952,n2949,n2951);
not gate_2933(n2953,n2952);
and gate_2934(n2954,n1839,n2953);
not gate_2935(n2955,n2954);
and gate_2936(n2956,n190,n522);
not gate_2937(n2957,n2956);
and gate_2938(n2958,pi9,n729);
and gate_2939(n2959,n1481,n2958);
not gate_2940(n2960,n2959);
and gate_2941(n2961,n2957,n2960);
not gate_2942(n2962,n2961);
and gate_2943(n2963,pi5,n2962);
not gate_2944(n2964,n2963);
and gate_2945(n2965,n25,n188);
and gate_2946(n2966,n1476,n2965);
not gate_2947(n2967,n2966);
and gate_2948(n2968,n2964,n2967);
not gate_2949(n2969,n2968);
and gate_2950(n2970,pi4,n2969);
not gate_2951(n2971,n2970);
and gate_2952(n2972,pi1,n25);
not gate_2953(n2973,n2972);
and gate_2954(n2974,pi1,n188);
not gate_2955(n2975,n2974);
and gate_2956(n2976,n322,n2975);
not gate_2957(n2977,n2976);
and gate_2958(n2978,n2973,n2977);
and gate_2959(n2979,n995,n2978);
not gate_2960(n2980,n2979);
and gate_2961(n2981,n2971,n2980);
not gate_2962(n2982,n2981);
and gate_2963(n2983,pi6,n2982);
not gate_2964(n2984,n2983);
and gate_2965(n2985,n1125,n1424);
and gate_2966(n2986,n306,n2985);
not gate_2967(n2987,n2986);
and gate_2968(n2988,n2984,n2987);
not gate_2969(n2989,n2988);
and gate_2970(n2990,pi0,n2989);
not gate_2971(n2991,n2990);
and gate_2972(n2992,n587,n1494);
not gate_2973(n2993,n2992);
and gate_2974(n2994,n26,n2993);
not gate_2975(n2995,n2994);
and gate_2976(n2996,n1217,n2995);
not gate_2977(n2997,n2996);
and gate_2978(n2998,n25,n2997);
not gate_2979(n2999,n2998);
and gate_2980(n3000,n234,n2533);
not gate_2981(n3001,n3000);
and gate_2982(n3002,n2999,n3001);
not gate_2983(n3003,n3002);
and gate_2984(n3004,n23,n3003);
not gate_2985(n3005,n3004);
and gate_2986(n3006,n21,n840);
and gate_2987(n3007,n1999,n3006);
not gate_2988(n3008,n3007);
and gate_2989(n3009,n3005,n3008);
not gate_2990(n3010,n3009);
and gate_2991(n3011,n1292,n3010);
not gate_2992(n3012,n3011);
and gate_2993(n3013,n2991,n3012);
and gate_2994(n3014,n2955,n3013);
not gate_2995(n3015,n3014);
and gate_2996(n3016,n22,n3015);
not gate_2997(n3017,n3016);
and gate_2998(n3018,n20,n1154);
not gate_2999(n3019,n3018);
and gate_3000(n3020,n1153,n3019);
not gate_3001(n3021,n3020);
and gate_3002(n3022,n27,n3021);
not gate_3003(n3023,n3022);
and gate_3004(n3024,pi0,pi7);
not gate_3005(n3025,n3024);
and gate_3006(n3026,n1236,n3024);
not gate_3007(n3027,n3026);
and gate_3008(n3028,n3023,n3027);
not gate_3009(n3029,n3028);
and gate_3010(n3030,pi3,n3029);
not gate_3011(n3031,n3030);
and gate_3012(n3032,n23,n1154);
and gate_3013(n3033,pi0,n3032);
not gate_3014(n3034,n3033);
and gate_3015(n3035,n3031,n3034);
not gate_3016(n3036,n3035);
and gate_3017(n3037,pi1,n3036);
not gate_3018(n3038,n3037);
and gate_3019(n3039,pi0,n1235);
and gate_3020(n3040,n1072,n3039);
not gate_3021(n3041,n3040);
and gate_3022(n3042,n159,n2433);
not gate_3023(n3043,n3042);
and gate_3024(n3044,n3041,n3043);
not gate_3025(n3045,n3044);
and gate_3026(n3046,pi7,n3045);
not gate_3027(n3047,n3046);
and gate_3028(n3048,n1206,n2761);
not gate_3029(n3049,n3048);
and gate_3030(n3050,n3047,n3049);
not gate_3031(n3051,n3050);
and gate_3032(n3052,n21,n3051);
not gate_3033(n3053,n3052);
and gate_3034(n3054,n3038,n3053);
not gate_3035(n3055,n3054);
and gate_3036(n3056,pi5,n3055);
not gate_3037(n3057,n3056);
and gate_3038(n3058,n1199,n1334);
and gate_3039(n3059,n3025,n3058);
and gate_3040(n3060,n23,n3059);
not gate_3041(n3061,n3060);
and gate_3042(n3062,n1334,n2089);
and gate_3043(n3063,n1200,n3062);
not gate_3044(n3064,n3063);
and gate_3045(n3065,n3061,n3064);
not gate_3046(n3066,n3065);
and gate_3047(n3067,pi4,n3066);
not gate_3048(n3068,n3067);
and gate_3049(n3069,pi0,n522);
and gate_3050(n3070,n24,n1320);
and gate_3051(n3071,n3069,n3070);
not gate_3052(n3072,n3071);
and gate_3053(n3073,n3068,n3072);
not gate_3054(n3074,n3073);
and gate_3055(n3075,n25,n3074);
not gate_3056(n3076,n3075);
and gate_3057(n3077,n3057,n3076);
not gate_3058(n3078,n3077);
and gate_3059(n3079,pi9,n3078);
not gate_3060(n3080,n3079);
and gate_3061(n3081,n47,n1609);
not gate_3062(n3082,n3081);
and gate_3063(n3083,n25,n1324);
and gate_3064(n3084,n55,n3083);
not gate_3065(n3085,n3084);
and gate_3066(n3086,n3082,n3085);
and gate_3067(n3087,n76,n2741);
not gate_3068(n3088,n3087);
and gate_3069(n3089,n350,n557);
not gate_3070(n3090,n3089);
and gate_3071(n3091,n3088,n3090);
not gate_3072(n3092,n3091);
and gate_3073(n3093,n24,n3092);
not gate_3074(n3094,n3093);
and gate_3075(n3095,n3086,n3094);
not gate_3076(n3096,n3095);
and gate_3077(n3097,pi3,n3096);
not gate_3078(n3098,n3097);
and gate_3079(n3099,n76,n106);
not gate_3080(n3100,n3099);
and gate_3081(n3101,n24,n1625);
not gate_3082(n3102,n3101);
and gate_3083(n3103,n1234,n3102);
not gate_3084(n3104,n3103);
and gate_3085(n3105,n84,n3104);
not gate_3086(n3106,n3105);
and gate_3087(n3107,n3100,n3106);
not gate_3088(n3108,n3107);
and gate_3089(n3109,pi7,n3108);
not gate_3090(n3110,n3109);
and gate_3091(n3111,n370,n1348);
and gate_3092(n3112,n20,n3111);
not gate_3093(n3113,n3112);
and gate_3094(n3114,n3110,n3113);
not gate_3095(n3115,n3114);
and gate_3096(n3116,n23,n3115);
not gate_3097(n3117,n3116);
and gate_3098(n3118,n3098,n3117);
not gate_3099(n3119,n3118);
and gate_3100(n3120,n29,n3119);
not gate_3101(n3121,n3120);
and gate_3102(n3122,n3080,n3121);
not gate_3103(n3123,n3122);
and gate_3104(n3124,pi2,n3123);
not gate_3105(n3125,n3124);
and gate_3106(n3126,n3017,n3125);
not gate_3107(n3127,n3126);
and gate_3108(n3128,pi8,n3127);
not gate_3109(n3129,n3128);
and gate_3110(n3130,pi0,n426);
not gate_3111(n3131,n3130);
and gate_3112(n3132,n20,n149);
not gate_3113(n3133,n3132);
and gate_3114(n3134,n3131,n3133);
not gate_3115(n3135,n3134);
and gate_3116(n3136,n23,n133);
not gate_3117(n3137,n3136);
and gate_3118(n3138,n1849,n3137);
not gate_3119(n3139,n3138);
and gate_3120(n3140,n3135,n3139);
not gate_3121(n3141,n3140);
and gate_3122(n3142,n256,n1492);
not gate_3123(n3143,n3142);
and gate_3124(n3144,pi6,n3143);
and gate_3125(n3145,n20,n3144);
not gate_3126(n3146,n3145);
and gate_3127(n3147,n1324,n1909);
not gate_3128(n3148,n3147);
and gate_3129(n3149,n3146,n3148);
not gate_3130(n3150,n3149);
and gate_3131(n3151,n949,n3150);
not gate_3132(n3152,n3151);
and gate_3133(n3153,n3141,n3152);
not gate_3134(n3154,n3153);
and gate_3135(n3155,pi1,n3154);
not gate_3136(n3156,n3155);
and gate_3137(n3157,pi7,n537);
and gate_3138(n3158,pi6,n3157);
not gate_3139(n3159,n3158);
and gate_3140(n3160,n2110,n3159);
not gate_3141(n3161,n3160);
and gate_3142(n3162,n182,n2109);
not gate_3143(n3163,n3162);
and gate_3144(n3164,n3161,n3163);
and gate_3145(n3165,pi3,n3164);
not gate_3146(n3166,n3165);
and gate_3147(n3167,n20,n842);
and gate_3148(n3168,n1293,n3167);
not gate_3149(n3169,n3168);
and gate_3150(n3170,n3166,n3169);
not gate_3151(n3171,n3170);
and gate_3152(n3172,n21,n3171);
not gate_3153(n3173,n3172);
and gate_3154(n3174,n3156,n3173);
not gate_3155(n3175,n3174);
and gate_3156(n3176,pi2,n3175);
not gate_3157(n3177,n3176);
and gate_3158(n3178,n1329,n2181);
not gate_3159(n3179,n3178);
and gate_3160(n3180,n3088,n3179);
not gate_3161(n3181,n3180);
and gate_3162(n3182,pi9,n3181);
not gate_3163(n3183,n3182);
and gate_3164(n3184,n20,n90);
not gate_3165(n3185,n3184);
and gate_3166(n3186,pi0,n26);
not gate_3167(n3187,n3186);
and gate_3168(n3188,n3185,n3187);
and gate_3169(n3189,n181,n3188);
and gate_3170(n3190,pi1,n3189);
not gate_3171(n3191,n3190);
and gate_3172(n3192,n3183,n3191);
not gate_3173(n3193,n3192);
and gate_3174(n3194,pi3,n3193);
not gate_3175(n3195,n3194);
and gate_3176(n3196,n76,n1989);
not gate_3177(n3197,n3196);
and gate_3178(n3198,n160,n1627);
and gate_3179(n3199,n909,n3198);
not gate_3180(n3200,n3199);
and gate_3181(n3201,n3197,n3200);
not gate_3182(n3202,n3201);
and gate_3183(n3203,n448,n3202);
not gate_3184(n3204,n3203);
and gate_3185(n3205,n3195,n3204);
not gate_3186(n3206,n3205);
and gate_3187(n3207,n22,n3206);
not gate_3188(n3208,n3207);
and gate_3189(n3209,n3177,n3208);
not gate_3190(n3210,n3209);
and gate_3191(n3211,pi4,n3210);
not gate_3192(n3212,n3211);
and gate_3193(n3213,pi2,n927);
not gate_3194(n3214,n3213);
and gate_3195(n3215,n22,n949);
not gate_3196(n3216,n3215);
and gate_3197(n3217,n3214,n3216);
not gate_3198(n3218,n3217);
and gate_3199(n3219,n27,n3218);
not gate_3200(n3220,n3219);
and gate_3201(n3221,n22,n876);
not gate_3202(n3222,n3221);
and gate_3203(n3223,n3220,n3222);
not gate_3204(n3224,n3223);
and gate_3205(n3225,n26,n3224);
not gate_3206(n3226,n3225);
and gate_3207(n3227,n889,n1586);
not gate_3208(n3228,n3227);
and gate_3209(n3229,n3226,n3228);
not gate_3210(n3230,n3229);
and gate_3211(n3231,n20,n3230);
not gate_3212(n3232,n3231);
and gate_3213(n3233,n676,n1393);
not gate_3214(n3234,n3233);
and gate_3215(n3235,n1860,n3234);
not gate_3216(n3236,n3235);
and gate_3217(n3237,n27,n3236);
not gate_3218(n3238,n3237);
and gate_3219(n3239,n26,n190);
and gate_3220(n3240,n917,n3239);
not gate_3221(n3241,n3240);
and gate_3222(n3242,n3238,n3241);
not gate_3223(n3243,n3242);
and gate_3224(n3244,pi0,n3243);
not gate_3225(n3245,n3244);
and gate_3226(n3246,n3232,n3245);
not gate_3227(n3247,n3246);
and gate_3228(n3248,pi1,n3247);
not gate_3229(n3249,n3248);
and gate_3230(n3250,pi2,n324);
not gate_3231(n3251,n3250);
and gate_3232(n3252,n426,n1174);
not gate_3233(n3253,n3252);
and gate_3234(n3254,n3251,n3253);
not gate_3235(n3255,n3254);
and gate_3236(n3256,pi6,n3255);
not gate_3237(n3257,n3256);
and gate_3238(n3258,n925,n3083);
not gate_3239(n3259,n3258);
and gate_3240(n3260,n3257,n3259);
not gate_3241(n3261,n3260);
and gate_3242(n3262,pi0,n3261);
not gate_3243(n3263,n3262);
and gate_3244(n3264,n20,n917);
and gate_3245(n3265,n1552,n3264);
not gate_3246(n3266,n3265);
and gate_3247(n3267,n3263,n3266);
not gate_3248(n3268,n3267);
and gate_3249(n3269,n21,n3268);
not gate_3250(n3270,n3269);
and gate_3251(n3271,n3249,n3270);
not gate_3252(n3272,n3271);
and gate_3253(n3273,n995,n3272);
not gate_3254(n3274,n3273);
and gate_3255(n3275,n3212,n3274);
not gate_3256(n3276,n3275);
and gate_3257(n3277,n28,n3276);
not gate_3258(n3278,n3277);
and gate_3259(n3279,n3129,n3278);
and gate_3260(n3280,n2947,n3279);
and gate_3261(n3281,n859,n1233);
and gate_3262(n3282,n20,n3281);
not gate_3263(n3283,n3282);
and gate_3264(n3284,pi0,n2430);
and gate_3265(n3285,n1125,n3284);
not gate_3266(n3286,n3285);
and gate_3267(n3287,n3283,n3286);
not gate_3268(n3288,n3287);
and gate_3269(n3289,n22,n3288);
not gate_3270(n3290,n3289);
and gate_3271(n3291,n1128,n1235);
and gate_3272(n3292,n30,n3291);
and gate_3273(n3293,pi0,n3292);
not gate_3274(n3294,n3293);
and gate_3275(n3295,n3290,n3294);
not gate_3276(n3296,n3295);
and gate_3277(n3297,pi8,n3296);
not gate_3278(n3298,n3297);
and gate_3279(n3299,n247,n1154);
and gate_3280(n3300,n2439,n3299);
not gate_3281(n3301,n3300);
and gate_3282(n3302,n3298,n3301);
not gate_3283(n3303,n3302);
and gate_3284(n3304,n1483,n3303);
and gate_3285(n3305,n223,n3304);
not gate_3286(n3306,n3305);
and gate_3287(n3307,n3280,n3306);
and gate_3288(n3308,n2919,n3307);
and gate_3289(n3309,n20,n995);
and gate_3290(n3310,n2920,n3309);
not gate_3291(n3311,n3310);
and gate_3292(n3312,n24,n424);
and gate_3293(n3313,pi0,n3312);
not gate_3294(n3314,n3313);
and gate_3295(n3315,n232,n1292);
not gate_3296(n3316,n3315);
and gate_3297(n3317,n3314,n3316);
not gate_3298(n3318,n3317);
and gate_3299(n3319,n1506,n3318);
not gate_3300(n3320,n3319);
and gate_3301(n3321,n3311,n3320);
not gate_3302(n3322,n3321);
and gate_3303(n3323,n21,n3322);
not gate_3304(n3324,n3323);
and gate_3305(n3325,pi0,n1476);
and gate_3306(n3326,n419,n1233);
and gate_3307(n3327,n3325,n3326);
not gate_3308(n3328,n3327);
and gate_3309(n3329,n3324,n3328);
not gate_3310(n3330,n3329);
and gate_3311(n3331,n924,n3330);
and gate_3312(n3332,n920,n3331);
not gate_3313(n3333,n3332);
and gate_3314(n3334,n3308,n3333);
and gate_3315(n3335,n21,n288);
and gate_3316(n3336,n1019,n1674);
and gate_3317(n3337,n3335,n3336);
not gate_3318(n3338,n3337);
and gate_3319(n3339,n80,n1781);
not gate_3320(n3340,n3339);
and gate_3321(n3341,n74,n2124);
not gate_3322(n3342,n3341);
and gate_3323(n3343,n3340,n3342);
not gate_3324(n3344,n3343);
and gate_3325(n3345,n945,n3344);
not gate_3326(n3346,n3345);
and gate_3327(n3347,n3338,n3346);
not gate_3328(n3348,n3347);
and gate_3329(n3349,n192,n3348);
and gate_3330(n3350,n1300,n3349);
not gate_3331(n3351,n3350);
and gate_3332(n3352,n3334,n3351);
not gate_3333(po5,n3352);
and gate_3334(n3354,n22,n2430);
and gate_3335(n3355,n2408,n3354);
not gate_3336(n3356,n3355);
and gate_3337(n3357,pi2,n1072);
not gate_3338(n3358,n3357);
and gate_3339(n3359,n356,n810);
and gate_3340(n3360,pi7,n3359);
and gate_3341(n3361,n3357,n3360);
not gate_3342(n3362,n3361);
and gate_3343(n3363,n3356,n3362);
not gate_3344(n3364,n3363);
and gate_3345(n3365,n26,n3364);
not gate_3346(n3366,n3365);
and gate_3347(n3367,n22,n1674);
and gate_3348(n3368,n222,n843);
and gate_3349(n3369,n24,n3368);
and gate_3350(n3370,n3367,n3369);
not gate_3351(n3371,n3370);
and gate_3352(n3372,n3366,n3371);
not gate_3353(n3373,n3372);
and gate_3354(n3374,n29,n3373);
not gate_3355(n3375,n3374);
and gate_3356(n3376,pi3,n32);
not gate_3357(n3377,n3376);
and gate_3358(n3378,n22,pi6);
not gate_3359(n3379,n3378);
and gate_3360(n3380,n1455,n3379);
not gate_3361(n3381,n3380);
and gate_3362(n3382,n223,n3381);
and gate_3363(n3383,pi4,n3382);
and gate_3364(n3384,n3376,n3383);
not gate_3365(n3385,n3384);
and gate_3366(n3386,n3375,n3385);
not gate_3367(n3387,n3386);
and gate_3368(n3388,n564,n3387);
not gate_3369(n3389,n3388);
and gate_3370(n3390,pi5,n179);
not gate_3371(n3391,n3390);
and gate_3372(n3392,n25,n181);
not gate_3373(n3393,n3392);
and gate_3374(n3394,n3391,n3393);
not gate_3375(n3395,n3394);
and gate_3376(n3396,n23,pi6);
and gate_3377(n3397,n76,n3396);
not gate_3378(n3398,n3397);
and gate_3379(n3399,n84,n1820);
not gate_3380(n3400,n3399);
and gate_3381(n3401,n3398,n3400);
not gate_3382(n3402,n3401);
and gate_3383(n3403,n3395,n3402);
not gate_3384(n3404,n3403);
and gate_3385(n3405,pi7,n1334);
not gate_3386(n3406,n3405);
and gate_3387(n3407,n20,n166);
not gate_3388(n3408,n3407);
and gate_3389(n3409,n3406,n3408);
not gate_3390(n3410,n3409);
and gate_3391(n3411,n583,n3410);
and gate_3392(n3412,n23,n3411);
not gate_3393(n3413,n3412);
and gate_3394(n3414,n1586,n3325);
not gate_3395(n3415,n3414);
and gate_3396(n3416,n3413,n3415);
not gate_3397(n3417,n3416);
and gate_3398(n3418,n25,n3417);
not gate_3399(n3419,n3418);
and gate_3400(n3420,n183,n587);
and gate_3401(n3421,n90,n3420);
and gate_3402(n3422,n2774,n3421);
not gate_3403(n3423,n3422);
and gate_3404(n3424,n3419,n3423);
and gate_3405(n3425,n3404,n3424);
not gate_3406(n3426,n3425);
and gate_3407(n3427,n24,n3426);
not gate_3408(n3428,n3427);
and gate_3409(n3429,n605,n1276);
not gate_3410(n3430,n3429);
and gate_3411(n3431,n586,n1839);
not gate_3412(n3432,n3431);
and gate_3413(n3433,n3430,n3432);
not gate_3414(n3434,n3433);
and gate_3415(n3435,n1300,n3434);
not gate_3416(n3436,n3435);
and gate_3417(n3437,pi0,n2495);
not gate_3418(n3438,n3437);
and gate_3419(n3439,n20,n1123);
not gate_3420(n3440,n3439);
and gate_3421(n3441,n3438,n3440);
not gate_3422(n3442,n3441);
and gate_3423(n3443,n23,n3442);
not gate_3424(n3444,n3443);
and gate_3425(n3445,n133,n531);
not gate_3426(n3446,n3445);
and gate_3427(n3447,n3444,n3446);
not gate_3428(n3448,n3447);
and gate_3429(n3449,n21,n3448);
not gate_3430(n3450,n3449);
and gate_3431(n3451,n76,n620);
not gate_3432(n3452,n3451);
and gate_3433(n3453,n3450,n3452);
not gate_3434(n3454,n3453);
and gate_3435(n3455,pi7,n3454);
not gate_3436(n3456,n3455);
and gate_3437(n3457,n84,n123);
not gate_3438(n3458,n3457);
and gate_3439(n3459,n76,n1128);
not gate_3440(n3460,n3459);
and gate_3441(n3461,n3458,n3460);
not gate_3442(n3462,n3461);
and gate_3443(n3463,n1491,n3462);
not gate_3444(n3464,n3463);
and gate_3445(n3465,n3456,n3464);
not gate_3446(n3466,n3465);
and gate_3447(n3467,pi5,n3466);
not gate_3448(n3468,n3467);
and gate_3449(n3469,n55,n1320);
not gate_3450(n3470,n3469);
and gate_3451(n3471,n47,n1324);
not gate_3452(n3472,n3471);
and gate_3453(n3473,n3470,n3472);
and gate_3454(n3474,n76,n2533);
not gate_3455(n3475,n3474);
and gate_3456(n3476,n3473,n3475);
not gate_3457(n3477,n3476);
and gate_3458(n3478,pi3,n3477);
not gate_3459(n3479,n3478);
and gate_3460(n3480,pi0,n945);
and gate_3461(n3481,n1293,n3480);
not gate_3462(n3482,n3481);
and gate_3463(n3483,n3479,n3482);
not gate_3464(n3484,n3483);
and gate_3465(n3485,n25,n3484);
not gate_3466(n3486,n3485);
and gate_3467(n3487,n3468,n3486);
and gate_3468(n3488,n3436,n3487);
not gate_3469(n3489,n3488);
and gate_3470(n3490,pi4,n3489);
not gate_3471(n3491,n3490);
and gate_3472(n3492,n3428,n3491);
not gate_3473(n3493,n3492);
and gate_3474(n3494,n22,n3493);
not gate_3475(n3495,n3494);
and gate_3476(n3496,n810,n2370);
and gate_3477(n3497,n48,n3496);
and gate_3478(n3498,n24,n3497);
not gate_3479(n3499,n3498);
and gate_3480(n3500,pi4,n2368);
not gate_3481(n3501,n3500);
and gate_3482(n3502,n3499,n3501);
not gate_3483(n3503,n3502);
and gate_3484(n3504,pi9,n3503);
not gate_3485(n3505,n3504);
and gate_3486(n3506,n1750,n3325);
not gate_3487(n3507,n3506);
and gate_3488(n3508,n3505,n3507);
not gate_3489(n3509,n3508);
and gate_3490(n3510,n1453,n3509);
not gate_3491(n3511,n3510);
and gate_3492(n3512,n21,n2631);
not gate_3493(n3513,n3512);
and gate_3494(n3514,n1324,n2972);
not gate_3495(n3515,n3514);
and gate_3496(n3516,n3513,n3515);
not gate_3497(n3517,n3516);
and gate_3498(n3518,n20,n3517);
not gate_3499(n3519,n3518);
and gate_3500(n3520,n1145,n1452);
and gate_3501(n3521,n163,n3520);
not gate_3502(n3522,n3521);
and gate_3503(n3523,n3519,n3522);
not gate_3504(n3524,n3523);
and gate_3505(n3525,pi3,n3524);
not gate_3506(n3526,n3525);
and gate_3507(n3527,n55,n1625);
not gate_3508(n3528,n3527);
and gate_3509(n3529,n47,n1393);
not gate_3510(n3530,n3529);
and gate_3511(n3531,n3528,n3530);
not gate_3512(n3532,n3531);
and gate_3513(n3533,pi7,n3532);
not gate_3514(n3534,n3533);
and gate_3515(n3535,n350,n3407);
not gate_3516(n3536,n3535);
and gate_3517(n3537,n3534,n3536);
not gate_3518(n3538,n3537);
and gate_3519(n3539,n23,n3538);
not gate_3520(n3540,n3539);
and gate_3521(n3541,n3526,n3540);
not gate_3522(n3542,n3541);
and gate_3523(n3543,pi4,n3542);
not gate_3524(n3544,n3543);
and gate_3525(n3545,n350,n1197);
not gate_3526(n3546,n3545);
and gate_3527(n3547,n166,n370);
not gate_3528(n3548,n3547);
and gate_3529(n3549,n3546,n3548);
not gate_3530(n3550,n3549);
and gate_3531(n3551,pi0,n3550);
not gate_3532(n3552,n3551);
and gate_3533(n3553,n1420,n1429);
not gate_3534(n3554,n3553);
and gate_3535(n3555,n25,n3554);
not gate_3536(n3556,n3555);
and gate_3537(n3557,n234,n1197);
not gate_3538(n3558,n3557);
and gate_3539(n3559,n3556,n3558);
not gate_3540(n3560,n3559);
and gate_3541(n3561,n20,n3560);
not gate_3542(n3562,n3561);
and gate_3543(n3563,n3552,n3562);
not gate_3544(n3564,n3563);
and gate_3545(n3565,n995,n3564);
not gate_3546(n3566,n3565);
and gate_3547(n3567,n3544,n3566);
not gate_3548(n3568,n3567);
and gate_3549(n3569,pi9,n3568);
not gate_3550(n3570,n3569);
and gate_3551(n3571,n76,n90);
not gate_3552(n3572,n3571);
and gate_3553(n3573,n2371,n3186);
not gate_3554(n3574,n3573);
and gate_3555(n3575,n3572,n3574);
not gate_3556(n3576,n3575);
and gate_3557(n3577,n24,n3576);
not gate_3558(n3578,n3577);
and gate_3559(n3579,n20,n1063);
not gate_3560(n3580,n3579);
and gate_3561(n3581,n3578,n3580);
not gate_3562(n3582,n3581);
and gate_3563(n3583,pi7,n3582);
not gate_3564(n3584,n3583);
and gate_3565(n3585,n20,n1335);
not gate_3566(n3586,n3585);
and gate_3567(n3587,pi0,n1419);
not gate_3568(n3588,n3587);
and gate_3569(n3589,n3586,n3588);
not gate_3570(n3590,n3589);
and gate_3571(n3591,n153,n3590);
and gate_3572(n3592,pi4,n3591);
not gate_3573(n3593,n3592);
and gate_3574(n3594,n3584,n3593);
not gate_3575(n3595,n3594);
and gate_3576(n3596,n23,n3595);
not gate_3577(n3597,n3596);
and gate_3578(n3598,n98,n153);
not gate_3579(n3599,n3598);
and gate_3580(n3600,n552,n1024);
not gate_3581(n3601,n3600);
and gate_3582(n3602,n3599,n3601);
not gate_3583(n3603,n3602);
and gate_3584(n3604,n1504,n3603);
and gate_3585(n3605,n20,n3604);
not gate_3586(n3606,n3605);
and gate_3587(n3607,n3597,n3606);
not gate_3588(n3608,n3607);
and gate_3589(n3609,n29,n3608);
not gate_3590(n3610,n3609);
and gate_3591(n3611,n3570,n3610);
and gate_3592(n3612,n3511,n3611);
not gate_3593(n3613,n3612);
and gate_3594(n3614,pi2,n3613);
not gate_3595(n3615,n3614);
and gate_3596(n3616,n3495,n3615);
not gate_3597(n3617,n3616);
and gate_3598(n3618,pi8,n3617);
not gate_3599(n3619,n3618);
and gate_3600(n3620,n1005,n1999);
not gate_3601(n3621,n3620);
and gate_3602(n3622,n1207,n2709);
not gate_3603(n3623,n3622);
and gate_3604(n3624,n586,n3623);
not gate_3605(n3625,n3624);
and gate_3606(n3626,n3621,n3625);
not gate_3607(n3627,n3626);
and gate_3608(n3628,n30,n3627);
and gate_3609(n3629,pi0,n3628);
not gate_3610(n3630,n3629);
and gate_3611(n3631,pi0,n1003);
and gate_3612(n3632,n1360,n3631);
not gate_3613(n3633,n3632);
and gate_3614(n3634,n1004,n1481);
and gate_3615(n3635,n1602,n3634);
and gate_3616(n3636,n159,n3635);
not gate_3617(n3637,n3636);
and gate_3618(n3638,n3633,n3637);
not gate_3619(n3639,n3638);
and gate_3620(n3640,n37,n3639);
not gate_3621(n3641,n3640);
and gate_3622(n3642,n3630,n3641);
and gate_3623(n3643,n892,n1554);
not gate_3624(n3644,n3643);
and gate_3625(n3645,n2552,n3644);
and gate_3626(n3646,pi0,n3645);
not gate_3627(n3647,n3646);
and gate_3628(n3648,n51,n68);
not gate_3629(n3649,n3648);
and gate_3630(n3650,n3647,n3649);
not gate_3631(n3651,n3650);
and gate_3632(n3652,pi6,n3651);
not gate_3633(n3653,n3652);
and gate_3634(n3654,n1197,n2371);
and gate_3635(n3655,n699,n3654);
not gate_3636(n3656,n3655);
and gate_3637(n3657,n3653,n3656);
and gate_3638(n3658,n338,n1098);
not gate_3639(n3659,n3658);
and gate_3640(n3660,n181,n3659);
not gate_3641(n3661,n3660);
and gate_3642(n3662,n68,n179);
not gate_3643(n3663,n3662);
and gate_3644(n3664,n3661,n3663);
not gate_3645(n3665,n3664);
and gate_3646(n3666,n25,n3665);
not gate_3647(n3667,n3666);
and gate_3648(n3668,n510,n3390);
not gate_3649(n3669,n3668);
and gate_3650(n3670,n3667,n3669);
not gate_3651(n3671,n3670);
and gate_3652(n3672,pi6,n3671);
not gate_3653(n3673,n3672);
and gate_3654(n3674,n56,n690);
not gate_3655(n3675,n3674);
and gate_3656(n3676,n363,n2181);
not gate_3657(n3677,n3676);
and gate_3658(n3678,n3675,n3677);
not gate_3659(n3679,n3678);
and gate_3660(n3680,n21,n3679);
not gate_3661(n3681,n3680);
and gate_3662(n3682,n76,n2583);
not gate_3663(n3683,n3682);
and gate_3664(n3684,n3681,n3683);
not gate_3665(n3685,n3684);
and gate_3666(n3686,n133,n3685);
not gate_3667(n3687,n3686);
and gate_3668(n3688,n3673,n3687);
not gate_3669(n3689,n3688);
and gate_3670(n3690,n24,n3689);
not gate_3671(n3691,n3690);
and gate_3672(n3692,n123,n1287);
not gate_3673(n3693,n3692);
and gate_3674(n3694,n133,n1097);
not gate_3675(n3695,n3694);
and gate_3676(n3696,n3693,n3695);
not gate_3677(n3697,n3696);
and gate_3678(n3698,n27,n3697);
not gate_3679(n3699,n3698);
and gate_3680(n3700,n538,n1335);
and gate_3681(n3701,n1115,n3700);
and gate_3682(n3702,pi7,n3701);
not gate_3683(n3703,n3702);
and gate_3684(n3704,n3699,n3703);
not gate_3685(n3705,n3704);
and gate_3686(n3706,pi5,n3705);
not gate_3687(n3707,n3706);
and gate_3688(n3708,n1331,n3472);
not gate_3689(n3709,n3708);
and gate_3690(n3710,n822,n3709);
and gate_3691(n3711,n22,n3710);
not gate_3692(n3712,n3711);
and gate_3693(n3713,n3707,n3712);
not gate_3694(n3714,n3713);
and gate_3695(n3715,pi4,n3714);
not gate_3696(n3716,n3715);
and gate_3697(n3717,n3691,n3716);
and gate_3698(n3718,n3657,n3717);
not gate_3699(n3719,n3718);
and gate_3700(n3720,n23,n3719);
not gate_3701(n3721,n3720);
and gate_3702(n3722,n52,n59);
not gate_3703(n3723,n3722);
and gate_3704(n3724,n681,n3723);
not gate_3705(n3725,n3724);
and gate_3706(n3726,pi4,n121);
and gate_3707(n3727,n712,n3726);
not gate_3708(n3728,n3727);
and gate_3709(n3729,n921,n2733);
not gate_3710(n3730,n3729);
and gate_3711(n3731,n3728,n3730);
not gate_3712(n3732,n3731);
and gate_3713(n3733,pi7,n3732);
not gate_3714(n3734,n3733);
and gate_3715(n3735,n385,n3674);
not gate_3716(n3736,n3735);
and gate_3717(n3737,n3734,n3736);
and gate_3718(n3738,n3725,n3737);
not gate_3719(n3739,n3738);
and gate_3720(n3740,pi6,n3739);
not gate_3721(n3741,n3740);
and gate_3722(n3742,n80,n2965);
not gate_3723(n3743,n3742);
and gate_3724(n3744,n74,n1599);
not gate_3725(n3745,n3744);
and gate_3726(n3746,n3743,n3745);
not gate_3727(n3747,n3746);
and gate_3728(n3748,n20,n3747);
not gate_3729(n3749,n3748);
and gate_3730(n3750,n361,n1423);
and gate_3731(n3751,n121,n3750);
and gate_3732(n3752,pi0,n3751);
not gate_3733(n3753,n3752);
and gate_3734(n3754,n3749,n3753);
not gate_3735(n3755,n3754);
and gate_3736(n3756,n26,n3755);
not gate_3737(n3757,n3756);
and gate_3738(n3758,n3741,n3757);
not gate_3739(n3759,n3758);
and gate_3740(n3760,pi1,n3759);
not gate_3741(n3761,n3760);
and gate_3742(n3762,pi2,n153);
not gate_3743(n3763,n3762);
and gate_3744(n3764,n889,n1320);
not gate_3745(n3765,n3764);
and gate_3746(n3766,n3763,n3765);
not gate_3747(n3767,n3766);
and gate_3748(n3768,n29,n3767);
not gate_3749(n3769,n3768);
and gate_3750(n3770,n889,n1293);
not gate_3751(n3771,n3770);
and gate_3752(n3772,n3769,n3771);
not gate_3753(n3773,n3772);
and gate_3754(n3774,pi0,n3773);
not gate_3755(n3775,n3774);
and gate_3756(n3776,n465,n1176);
and gate_3757(n3777,n3379,n3776);
and gate_3758(n3778,n1336,n3777);
not gate_3759(n3779,n3778);
and gate_3760(n3780,n3775,n3779);
not gate_3761(n3781,n3780);
and gate_3762(n3782,n24,n3781);
not gate_3763(n3783,n3782);
and gate_3764(n3784,pi2,n3395);
not gate_3765(n3785,n3784);
and gate_3766(n3786,n131,n190);
not gate_3767(n3787,n3786);
and gate_3768(n3788,n3785,n3787);
not gate_3769(n3789,n3788);
and gate_3770(n3790,n26,n3789);
not gate_3771(n3791,n3790);
and gate_3772(n3792,n131,n1999);
not gate_3773(n3793,n3792);
and gate_3774(n3794,n3791,n3793);
not gate_3775(n3795,n3794);
and gate_3776(n3796,n1292,n3795);
not gate_3777(n3797,n3796);
and gate_3778(n3798,n3783,n3797);
not gate_3779(n3799,n3798);
and gate_3780(n3800,n21,n3799);
not gate_3781(n3801,n3800);
and gate_3782(n3802,n3761,n3801);
not gate_3783(n3803,n3802);
and gate_3784(n3804,pi3,n3803);
not gate_3785(n3805,n3804);
and gate_3786(n3806,n3721,n3805);
and gate_3787(n3807,n3642,n3806);
not gate_3788(n3808,n3807);
and gate_3789(n3809,n28,n3808);
not gate_3790(n3810,n3809);
and gate_3791(n3811,n3619,n3810);
and gate_3792(n3812,n3389,n3811);
not gate_3793(po6,n3812);
and gate_3794(n3814,n55,n1686);
not gate_3795(n3815,n3814);
and gate_3796(n3816,n570,n1292);
not gate_3797(n3817,n3816);
and gate_3798(n3818,n3815,n3817);
not gate_3799(n3819,n3818);
and gate_3800(n3820,n25,n3819);
not gate_3801(n3821,n3820);
and gate_3802(n3822,n24,n211);
and gate_3803(n3823,n47,n3822);
not gate_3804(n3824,n3823);
and gate_3805(n3825,n3821,n3824);
not gate_3806(n3826,n3825);
and gate_3807(n3827,n1452,n1508);
and gate_3808(n3828,n2495,n3827);
and gate_3809(n3829,n3826,n3828);
not gate_3810(n3830,n3829);
and gate_3811(n3831,pi1,n1809);
not gate_3812(n3832,n3831);
and gate_3813(n3833,n1179,n3832);
not gate_3814(n3834,n3833);
and gate_3815(n3835,pi5,n3834);
not gate_3816(n3836,n3835);
and gate_3817(n3837,n203,n1005);
not gate_3818(n3838,n3837);
and gate_3819(n3839,n3836,n3838);
not gate_3820(n3840,n3839);
and gate_3821(n3841,pi0,n3840);
not gate_3822(n3842,n3841);
and gate_3823(n3843,n21,n208);
not gate_3824(n3844,n3843);
and gate_3825(n3845,pi1,n211);
not gate_3826(n3846,n3845);
and gate_3827(n3847,n3844,n3846);
not gate_3828(n3848,n3847);
and gate_3829(n3849,n1292,n3848);
not gate_3830(n3850,n3849);
and gate_3831(n3851,n3842,n3850);
not gate_3832(n3852,n3851);
and gate_3833(n3853,n29,n3852);
not gate_3834(n3854,n3853);
and gate_3835(n3855,pi0,n1690);
not gate_3836(n3856,n3855);
and gate_3837(n3857,n2734,n3856);
not gate_3838(n3858,n3857);
and gate_3839(n3859,n832,n3858);
and gate_3840(n3860,pi1,n3859);
not gate_3841(n3861,n3860);
and gate_3842(n3862,n3854,n3861);
not gate_3843(n3863,n3862);
and gate_3844(n3864,n23,n3863);
not gate_3845(n3865,n3864);
and gate_3846(n3866,n583,n2164);
not gate_3847(n3867,n3866);
and gate_3848(n3868,n21,n832);
not gate_3849(n3869,n3868);
and gate_3850(n3870,n3867,n3869);
not gate_3851(n3871,n3870);
and gate_3852(n3872,n28,n3871);
not gate_3853(n3873,n3872);
and gate_3854(n3874,n25,n278);
and gate_3855(n3875,n47,n3874);
not gate_3856(n3876,n3875);
and gate_3857(n3877,n3873,n3876);
not gate_3858(n3878,n3877);
and gate_3859(n3879,pi4,n3878);
not gate_3860(n3880,n3879);
and gate_3861(n3881,n442,n1005);
and gate_3862(n3882,n20,n3881);
not gate_3863(n3883,n3882);
and gate_3864(n3884,n3880,n3883);
not gate_3865(n3885,n3884);
and gate_3866(n3886,pi3,n3885);
not gate_3867(n3887,n3886);
and gate_3868(n3888,n3865,n3887);
not gate_3869(n3889,n3888);
and gate_3870(n3890,pi6,n3889);
not gate_3871(n3891,n3890);
and gate_3872(n3892,n76,n352);
not gate_3873(n3893,n3892);
and gate_3874(n3894,n84,n354);
not gate_3875(n3895,n3894);
and gate_3876(n3896,n3893,n3895);
and gate_3877(n3897,n2094,n2100);
and gate_3878(n3898,n564,n3897);
and gate_3879(n3899,n23,n3898);
not gate_3880(n3900,n3899);
and gate_3881(n3901,n3896,n3900);
not gate_3882(n3902,n3901);
and gate_3883(n3903,pi9,n3902);
not gate_3884(n3904,n3903);
and gate_3885(n3905,n20,n28);
not gate_3886(n3906,n3905);
and gate_3887(n3907,n329,n3906);
and gate_3888(n3908,n949,n3907);
and gate_3889(n3909,pi1,n3908);
not gate_3890(n3910,n3909);
and gate_3891(n3911,n3904,n3910);
not gate_3892(n3912,n3911);
and gate_3893(n3913,pi4,n3912);
not gate_3894(n3914,n3913);
and gate_3895(n3915,n278,n1019);
and gate_3896(n3916,n1905,n3915);
not gate_3897(n3917,n3916);
and gate_3898(n3918,n3914,n3917);
not gate_3899(n3919,n3918);
and gate_3900(n3920,n26,n3919);
not gate_3901(n3921,n3920);
and gate_3902(n3922,n3891,n3921);
not gate_3903(n3923,n3922);
and gate_3904(n3924,pi7,n3923);
not gate_3905(n3925,n3924);
and gate_3906(n3926,pi1,n771);
not gate_3907(n3927,n3926);
and gate_3908(n3928,n522,n766);
not gate_3909(n3929,n3928);
and gate_3910(n3930,n3927,n3929);
not gate_3911(n3931,n3930);
and gate_3912(n3932,pi8,n3931);
not gate_3913(n3933,n3932);
and gate_3914(n3934,n767,n2432);
and gate_3915(n3935,n567,n3934);
not gate_3916(n3936,n3935);
and gate_3917(n3937,n3933,n3936);
not gate_3918(n3938,n3937);
and gate_3919(n3939,pi0,n3938);
not gate_3920(n3940,n3939);
and gate_3921(n3941,n297,n3377);
not gate_3922(n3942,n3941);
and gate_3923(n3943,n21,n3942);
not gate_3924(n3944,n3943);
and gate_3925(n3945,n39,n1476);
not gate_3926(n3946,n3945);
and gate_3927(n3947,n3944,n3946);
not gate_3928(n3948,n3947);
and gate_3929(n3949,pi4,n3948);
not gate_3930(n3950,n3949);
and gate_3931(n3951,n522,n714);
not gate_3932(n3952,n3951);
and gate_3933(n3953,n3950,n3952);
not gate_3934(n3954,n3953);
and gate_3935(n3955,n20,n3954);
not gate_3936(n3956,n3955);
and gate_3937(n3957,n3940,n3956);
not gate_3938(n3958,n3957);
and gate_3939(n3959,n26,n3958);
not gate_3940(n3960,n3959);
and gate_3941(n3961,pi0,n605);
and gate_3942(n3962,n24,n39);
and gate_3943(n3963,n3961,n3962);
not gate_3944(n3964,n3963);
and gate_3945(n3965,n21,n39);
not gate_3946(n3966,n3965);
and gate_3947(n3967,pi3,n462);
not gate_3948(n3968,n3967);
and gate_3949(n3969,pi1,n3967);
not gate_3950(n3970,n3969);
and gate_3951(n3971,n3966,n3970);
not gate_3952(n3972,n3971);
and gate_3953(n3973,n1292,n3972);
not gate_3954(n3974,n3973);
and gate_3955(n3975,n3964,n3974);
not gate_3956(n3976,n3975);
and gate_3957(n3977,pi6,n3976);
not gate_3958(n3978,n3977);
and gate_3959(n3979,n3960,n3978);
not gate_3960(n3980,n3979);
and gate_3961(n3981,n25,n3980);
not gate_3962(n3982,n3981);
and gate_3963(n3983,n461,n582);
and gate_3964(n3984,n1145,n3983);
and gate_3965(n3985,n23,n3984);
not gate_3966(n3986,n3985);
and gate_3967(n3987,n26,n247);
and gate_3968(n3988,n522,n3987);
not gate_3969(n3989,n3988);
and gate_3970(n3990,n3986,n3989);
not gate_3971(n3991,n3990);
and gate_3972(n3992,pi0,n3991);
not gate_3973(n3993,n3992);
and gate_3974(n3994,n522,n1123);
not gate_3975(n3995,n3994);
and gate_3976(n3996,pi1,n1504);
not gate_3977(n3997,n3996);
and gate_3978(n3998,n1507,n3997);
not gate_3979(n3999,n3998);
and gate_3980(n4000,pi9,n3999);
not gate_3981(n4001,n4000);
and gate_3982(n4002,n3995,n4001);
not gate_3983(n4003,n4002);
and gate_3984(n4004,pi8,n4003);
not gate_3985(n4005,n4004);
and gate_3986(n4006,n1476,n3987);
not gate_3987(n4007,n4006);
and gate_3988(n4008,n4005,n4007);
not gate_3989(n4009,n4008);
and gate_3990(n4010,n20,n4009);
not gate_3991(n4011,n4010);
and gate_3992(n4012,n3993,n4011);
not gate_3993(n4013,n4012);
and gate_3994(n4014,n979,n4013);
not gate_3995(n4015,n4014);
and gate_3996(n4016,n3982,n4015);
not gate_3997(n4017,n4016);
and gate_3998(n4018,n27,n4017);
not gate_3999(n4019,n4018);
and gate_4000(n4020,n3925,n4019);
and gate_4001(n4021,n3830,n4020);
not gate_4002(n4022,n4021);
and gate_4003(n4023,pi2,n4022);
not gate_4004(n4024,n4023);
and gate_4005(n4025,n21,n1506);
not gate_4006(n4026,n4025);
and gate_4007(n4027,n3997,n4026);
not gate_4008(n4028,n4027);
and gate_4009(n4029,n121,n4028);
and gate_4010(n4030,n20,n4029);
not gate_4011(n4031,n4030);
and gate_4012(n4032,n125,n3325);
not gate_4013(n4033,n4032);
and gate_4014(n4034,n4031,n4033);
not gate_4015(n4035,n4034);
and gate_4016(n4036,n556,n4035);
not gate_4017(n4037,n4036);
and gate_4018(n4038,n729,n1299);
and gate_4019(n4039,n963,n4038);
and gate_4020(n4040,n25,n4039);
not gate_4021(n4041,n4040);
and gate_4022(n4042,pi9,n3143);
and gate_4023(n4043,n20,n4042);
not gate_4024(n4044,n4043);
and gate_4025(n4045,n114,n730);
not gate_4026(n4046,n4045);
and gate_4027(n4047,n4044,n4046);
not gate_4028(n4048,n4047);
and gate_4029(n4049,pi5,n4048);
not gate_4030(n4050,n4049);
and gate_4031(n4051,n4041,n4050);
not gate_4032(n4052,n4051);
and gate_4033(n4053,pi6,n4052);
not gate_4034(n4054,n4053);
and gate_4035(n4055,n1337,n3025);
not gate_4036(n4056,n4055);
and gate_4037(n4057,n2450,n4056);
and gate_4038(n4058,n69,n4057);
not gate_4039(n4059,n4058);
and gate_4040(n4060,n4054,n4059);
not gate_4041(n4061,n4060);
and gate_4042(n4062,n28,n4061);
not gate_4043(n4063,n4062);
and gate_4044(n4064,pi0,n1644);
not gate_4045(n4065,n4064);
and gate_4046(n4066,n1128,n2761);
not gate_4047(n4067,n4066);
and gate_4048(n4068,n4065,n4067);
not gate_4049(n4069,n4068);
and gate_4050(n4070,n153,n4069);
not gate_4051(n4071,n4070);
and gate_4052(n4072,n1609,n2774);
not gate_4053(n4073,n4072);
and gate_4054(n4074,n4071,n4073);
not gate_4055(n4075,n4074);
and gate_4056(n4076,pi8,n4075);
not gate_4057(n4077,n4076);
and gate_4058(n4078,n4063,n4077);
not gate_4059(n4079,n4078);
and gate_4060(n4080,n21,n4079);
not gate_4061(n4081,n4080);
and gate_4062(n4082,n829,n2831);
not gate_4063(n4083,n4082);
and gate_4064(n4084,n842,n2617);
not gate_4065(n4085,n4084);
and gate_4066(n4086,n4083,n4085);
not gate_4067(n4087,n4086);
and gate_4068(n4088,pi0,n4087);
not gate_4069(n4089,n4088);
and gate_4070(n4090,n858,n3144);
not gate_4071(n4091,n4090);
and gate_4072(n4092,n193,n1820);
not gate_4073(n4093,n4092);
and gate_4074(n4094,n4091,n4093);
not gate_4075(n4095,n4094);
and gate_4076(n4096,n2092,n4095);
and gate_4077(n4097,n20,n4096);
not gate_4078(n4098,n4097);
and gate_4079(n4099,n4089,n4098);
not gate_4080(n4100,n4099);
and gate_4081(n4101,pi1,n4100);
not gate_4082(n4102,n4101);
and gate_4083(n4103,n4081,n4102);
and gate_4084(n4104,n4037,n4103);
not gate_4085(n4105,n4104);
and gate_4086(n4106,pi4,n4105);
not gate_4087(n4107,n4106);
and gate_4088(n4108,n25,n421);
and gate_4089(n4109,n522,n4108);
not gate_4090(n4110,n4109);
and gate_4091(n4111,pi7,n357);
and gate_4092(n4112,n1025,n4111);
not gate_4093(n4113,n4112);
and gate_4094(n4114,n4110,n4113);
not gate_4095(n4115,n4114);
and gate_4096(n4116,n20,n4115);
not gate_4097(n4117,n4116);
and gate_4098(n4118,n25,n419);
and gate_4099(n4119,n3961,n4118);
not gate_4100(n4120,n4119);
and gate_4101(n4121,n4117,n4120);
not gate_4102(n4122,n4121);
and gate_4103(n4123,n1128,n4122);
not gate_4104(n4124,n4123);
and gate_4105(n4125,n232,n522);
not gate_4106(n4126,n4125);
and gate_4107(n4127,n565,n3143);
not gate_4108(n4128,n4127);
and gate_4109(n4129,n4126,n4128);
not gate_4110(n4130,n4129);
and gate_4111(n4131,n26,n4130);
not gate_4112(n4132,n4131);
and gate_4113(n4133,n522,n2182);
not gate_4114(n4134,n4133);
and gate_4115(n4135,n4132,n4134);
not gate_4116(n4136,n4135);
and gate_4117(n4137,pi9,n4136);
not gate_4118(n4138,n4137);
and gate_4119(n4139,n21,n372);
not gate_4120(n4140,n4139);
and gate_4121(n4141,n2245,n4140);
not gate_4122(n4142,n4141);
and gate_4123(n4143,pi6,n4142);
not gate_4124(n4144,n4143);
and gate_4125(n4145,n232,n1332);
not gate_4126(n4146,n4145);
and gate_4127(n4147,n4144,n4146);
not gate_4128(n4148,n4147);
and gate_4129(n4149,n960,n4148);
not gate_4130(n4150,n4149);
and gate_4131(n4151,n4138,n4150);
not gate_4132(n4152,n4151);
and gate_4133(n4153,n20,n4152);
not gate_4134(n4154,n4153);
and gate_4135(n4155,n26,n571);
not gate_4136(n4156,n4155);
and gate_4137(n4157,n194,n1483);
and gate_4138(n4158,n1128,n4157);
not gate_4139(n4159,n4158);
and gate_4140(n4160,n4156,n4159);
not gate_4141(n4161,n4160);
and gate_4142(n4162,n23,n4161);
not gate_4143(n4163,n4162);
and gate_4144(n4164,n278,n1320);
not gate_4145(n4165,n4164);
and gate_4146(n4166,n462,n1324);
not gate_4147(n4167,n4166);
and gate_4148(n4168,n4165,n4167);
not gate_4149(n4169,n4168);
and gate_4150(n4170,n1476,n4169);
not gate_4151(n4171,n4170);
and gate_4152(n4172,n4163,n4171);
not gate_4153(n4173,n4172);
and gate_4154(n4174,pi0,n4173);
not gate_4155(n4175,n4174);
and gate_4156(n4176,n4154,n4175);
not gate_4157(n4177,n4176);
and gate_4158(n4178,pi5,n4177);
not gate_4159(n4179,n4178);
and gate_4160(n4180,n20,n3139);
not gate_4161(n4181,n4180);
and gate_4162(n4182,n2774,n3239);
not gate_4163(n4183,n4182);
and gate_4164(n4184,n4181,n4183);
not gate_4165(n4185,n4184);
and gate_4166(n4186,n28,n4185);
not gate_4167(n4187,n4186);
and gate_4168(n4188,n1909,n2617);
not gate_4169(n4189,n4188);
and gate_4170(n4190,n4187,n4189);
not gate_4171(n4191,n4190);
and gate_4172(n4192,pi1,n4191);
not gate_4173(n4193,n4192);
and gate_4174(n4194,n281,n3968);
not gate_4175(n4195,n4194);
and gate_4176(n4196,n1352,n4195);
and gate_4177(n4197,pi0,n4196);
not gate_4178(n4198,n4197);
and gate_4179(n4199,n4193,n4198);
not gate_4180(n4200,n4199);
and gate_4181(n4201,n25,n4200);
not gate_4182(n4202,n4201);
and gate_4183(n4203,n4179,n4202);
and gate_4184(n4204,n4124,n4203);
not gate_4185(n4205,n4204);
and gate_4186(n4206,n24,n4205);
not gate_4187(n4207,n4206);
and gate_4188(n4208,n4107,n4207);
not gate_4189(n4209,n4208);
and gate_4190(n4210,n22,n4209);
not gate_4191(n4211,n4210);
and gate_4192(n4212,n4024,n4211);
not gate_4193(po7,n4212);
and gate_4194(n4214,n632,n3069);
not gate_4195(n4215,n4214);
and gate_4196(n4216,n3893,n4215);
not gate_4197(n4217,n4216);
and gate_4198(n4218,n466,n4217);
and gate_4199(n4219,n29,n4218);
not gate_4200(n4220,n4219);
and gate_4201(n4221,n32,n264);
and gate_4202(n4222,n1097,n4221);
not gate_4203(n4223,n4222);
and gate_4204(n4224,n4220,n4223);
not gate_4205(n4225,n4224);
and gate_4206(n4226,n24,n4225);
not gate_4207(n4227,n4226);
and gate_4208(n4228,n787,n3874);
and gate_4209(n4229,n20,n4228);
not gate_4210(n4230,n4229);
and gate_4211(n4231,n4227,n4230);
not gate_4212(n4232,n4231);
and gate_4213(n4233,n1453,n4232);
not gate_4214(n4234,n4233);
and gate_4215(n4235,n633,n810);
and gate_4216(n4236,n3143,n4235);
not gate_4217(n4237,n4236);
and gate_4218(n4238,n874,n2593);
not gate_4219(n4239,n4238);
and gate_4220(n4240,n4237,n4239);
not gate_4221(n4241,n4240);
and gate_4222(n4242,pi0,n4241);
not gate_4223(n4243,n4242);
and gate_4224(n4244,n463,n3143);
not gate_4225(n4245,n4244);
and gate_4226(n4246,n131,n730);
not gate_4227(n4247,n4246);
and gate_4228(n4248,n4245,n4247);
not gate_4229(n4249,n4248);
and gate_4230(n4250,pi8,n4249);
not gate_4231(n4251,n4250);
and gate_4232(n4252,n425,n920);
and gate_4233(n4253,n354,n4252);
not gate_4234(n4254,n4253);
and gate_4235(n4255,n4251,n4254);
not gate_4236(n4256,n4255);
and gate_4237(n4257,n20,n4256);
not gate_4238(n4258,n4257);
and gate_4239(n4259,n4243,n4258);
not gate_4240(n4260,n4259);
and gate_4241(n4261,pi4,n4260);
not gate_4242(n4262,n4261);
and gate_4243(n4263,pi8,n4056);
not gate_4244(n4264,n4263);
and gate_4245(n4265,n419,n990);
not gate_4246(n4266,n4265);
and gate_4247(n4267,n4264,n4266);
not gate_4248(n4268,n4267);
and gate_4249(n4269,pi5,n4268);
not gate_4250(n4270,n4269);
and gate_4251(n4271,n2391,n2393);
not gate_4252(n4272,n4271);
and gate_4253(n4273,n49,n4272);
not gate_4254(n4274,n4273);
and gate_4255(n4275,n4270,n4274);
not gate_4256(n4276,n4275);
and gate_4257(n4277,pi3,n4276);
not gate_4258(n4278,n4277);
and gate_4259(n4279,n163,n2896);
not gate_4260(n4280,n4279);
and gate_4261(n4281,n4278,n4280);
not gate_4262(n4282,n4281);
and gate_4263(n4283,n24,n4282);
not gate_4264(n4284,n4283);
and gate_4265(n4285,n4262,n4284);
not gate_4266(n4286,n4285);
and gate_4267(n4287,n21,n4286);
not gate_4268(n4288,n4287);
and gate_4269(n4289,n81,n1687);
not gate_4270(n4290,n4289);
and gate_4271(n4291,pi0,n24);
not gate_4272(n4292,n4291);
and gate_4273(n4293,n637,n4292);
not gate_4274(n4294,n4293);
and gate_4275(n4295,n4290,n4293);
not gate_4276(n4296,n4295);
and gate_4277(n4297,n4289,n4294);
not gate_4278(n4298,n4297);
and gate_4279(n4299,n4296,n4298);
not gate_4280(n4300,n4299);
and gate_4281(n4301,n27,n4300);
not gate_4282(n4302,n4301);
and gate_4283(n4303,pi0,pi8);
not gate_4284(n4304,n4303);
and gate_4285(n4305,n3906,n4304);
not gate_4286(n4306,n4305);
and gate_4287(n4307,n688,n4306);
and gate_4288(n4308,n22,n4307);
not gate_4289(n4309,n4308);
and gate_4290(n4310,n4302,n4309);
not gate_4291(n4311,n4310);
and gate_4292(n4312,pi3,n4311);
not gate_4293(n4313,n4312);
and gate_4294(n4314,n232,n2733);
not gate_4295(n4315,n4314);
and gate_4296(n4316,pi7,n1708);
and gate_4297(n4317,n2734,n4316);
not gate_4298(n4318,n4317);
and gate_4299(n4319,n4315,n4318);
not gate_4300(n4320,n4319);
and gate_4301(n4321,n37,n4320);
not gate_4302(n4322,n4321);
and gate_4303(n4323,n4313,n4322);
not gate_4304(n4324,n4323);
and gate_4305(n4325,pi5,n4324);
not gate_4306(n4326,n4325);
and gate_4307(n4327,pi3,n1709);
not gate_4308(n4328,n4327);
and gate_4309(n4329,n874,n1686);
not gate_4310(n4330,n4329);
and gate_4311(n4331,n4328,n4330);
not gate_4312(n4332,n4331);
and gate_4313(n4333,pi7,n4332);
not gate_4314(n4334,n4333);
and gate_4315(n4335,pi4,n2896);
not gate_4316(n4336,n4335);
and gate_4317(n4337,n4334,n4336);
not gate_4318(n4338,n4337);
and gate_4319(n4339,pi0,n4338);
not gate_4320(n4340,n4339);
and gate_4321(n4341,n24,n421);
and gate_4322(n4342,n2471,n4341);
not gate_4323(n4343,n4342);
and gate_4324(n4344,n4340,n4343);
not gate_4325(n4345,n4344);
and gate_4326(n4346,n25,n4345);
not gate_4327(n4347,n4346);
and gate_4328(n4348,n4326,n4347);
not gate_4329(n4349,n4348);
and gate_4330(n4350,pi1,n4349);
not gate_4331(n4351,n4350);
and gate_4332(n4352,n4288,n4351);
not gate_4333(n4353,n4352);
and gate_4334(n4354,pi9,n4353);
not gate_4335(n4355,n4354);
and gate_4336(n4356,pi0,n1178);
and gate_4337(n4357,n4118,n4356);
not gate_4338(n4358,n4357);
and gate_4339(n4359,n2081,n2733);
not gate_4340(n4360,n4359);
and gate_4341(n4361,n4358,n4360);
not gate_4342(n4362,n4361);
and gate_4343(n4363,n365,n4362);
not gate_4344(n4364,n4363);
and gate_4345(n4365,pi2,n845);
not gate_4346(n4366,n4365);
and gate_4347(n4367,n2379,n4366);
not gate_4348(n4368,n4367);
and gate_4349(n4369,n28,n4368);
not gate_4350(n4370,n4369);
and gate_4351(n4371,n37,n2092);
not gate_4352(n4372,n4371);
and gate_4353(n4373,n4370,n4372);
not gate_4354(n4374,n4373);
and gate_4355(n4375,n24,n4374);
not gate_4356(n4376,n4375);
and gate_4357(n4377,n613,n2093);
and gate_4358(n4378,n2430,n4377);
not gate_4359(n4379,n4378);
and gate_4360(n4380,n4376,n4379);
not gate_4361(n4381,n4380);
and gate_4362(n4382,pi1,n4381);
not gate_4363(n4383,n4382);
and gate_4364(n4384,n74,n2092);
not gate_4365(n4385,n4384);
and gate_4366(n4386,n612,n1058);
not gate_4367(n4387,n4386);
and gate_4368(n4388,n4385,n4387);
not gate_4369(n4389,n4388);
and gate_4370(n4390,n522,n4389);
not gate_4371(n4391,n4390);
and gate_4372(n4392,n4383,n4391);
not gate_4373(n4393,n4392);
and gate_4374(n4394,pi7,n4393);
not gate_4375(n4395,n4394);
and gate_4376(n4396,n810,n1071);
and gate_4377(n4397,n330,n4396);
and gate_4378(n4398,pi2,n4397);
not gate_4379(n4399,n4398);
and gate_4380(n4400,n205,n1648);
not gate_4381(n4401,n4400);
and gate_4382(n4402,n4399,n4401);
not gate_4383(n4403,n4402);
and gate_4384(n4404,n1480,n4403);
not gate_4385(n4405,n4404);
and gate_4386(n4406,n4395,n4405);
not gate_4387(n4407,n4406);
and gate_4388(n4408,pi0,n4407);
not gate_4389(n4409,n4408);
and gate_4390(n4410,n1071,n3831);
not gate_4391(n4411,n4410);
and gate_4392(n4412,n21,n356);
and gate_4393(n4413,n1809,n4412);
not gate_4394(n4414,n4413);
and gate_4395(n4415,n4411,n4414);
not gate_4396(n4416,n4415);
and gate_4397(n4417,pi7,n4416);
not gate_4398(n4418,n4417);
and gate_4399(n4419,n24,n4125);
not gate_4400(n4420,n4419);
and gate_4401(n4421,n4418,n4420);
not gate_4402(n4422,n4421);
and gate_4403(n4423,pi5,n4422);
not gate_4404(n4424,n4423);
and gate_4405(n4425,n1178,n4108);
not gate_4406(n4426,n4425);
and gate_4407(n4427,n4424,n4426);
not gate_4408(n4428,n4427);
and gate_4409(n4429,n22,n4428);
not gate_4410(n4430,n4429);
and gate_4411(n4431,n997,n4118);
not gate_4412(n4432,n4431);
and gate_4413(n4433,n1423,n1691);
and gate_4414(n4434,n1020,n4433);
and gate_4415(n4435,n605,n4434);
not gate_4416(n4436,n4435);
and gate_4417(n4437,n4432,n4436);
not gate_4418(n4438,n4437);
and gate_4419(n4439,pi2,n4438);
not gate_4420(n4440,n4439);
and gate_4421(n4441,n4430,n4440);
not gate_4422(n4442,n4441);
and gate_4423(n4443,n20,n4442);
not gate_4424(n4444,n4443);
and gate_4425(n4445,n4409,n4444);
and gate_4426(n4446,n4364,n4445);
not gate_4427(n4447,n4446);
and gate_4428(n4448,n29,n4447);
not gate_4429(n4449,n4448);
and gate_4430(n4450,n4355,n4449);
not gate_4431(n4451,n4450);
and gate_4432(n4452,n26,n4451);
not gate_4433(n4453,n4452);
and gate_4434(n4454,n810,n890);
and gate_4435(n4455,n181,n4454);
not gate_4436(n4456,n4455);
and gate_4437(n4457,n3222,n4456);
not gate_4438(n4458,n4457);
and gate_4439(n4459,n21,n4458);
not gate_4440(n4460,n4459);
and gate_4441(n4461,pi1,n288);
and gate_4442(n4462,n319,n4461);
not gate_4443(n4463,n4462);
and gate_4444(n4464,n4460,n4463);
not gate_4445(n4465,n4464);
and gate_4446(n4466,n20,n4465);
not gate_4447(n4467,n4466);
and gate_4448(n4468,n188,n304);
and gate_4449(n4469,n1070,n4468);
not gate_4450(n4470,n4469);
and gate_4451(n4471,n4467,n4470);
not gate_4452(n4472,n4471);
and gate_4453(n4473,n1809,n4472);
not gate_4454(n4474,n4473);
and gate_4455(n4475,n189,n4305);
not gate_4456(n4476,n4475);
and gate_4457(n4477,n191,n2097);
not gate_4458(n4478,n4477);
and gate_4459(n4479,n4476,n4478);
and gate_4460(n4480,n2433,n4479);
not gate_4461(n4481,n4480);
and gate_4462(n4482,n267,n3284);
not gate_4463(n4483,n4482);
and gate_4464(n4484,n4481,n4483);
not gate_4465(n4485,n4484);
and gate_4466(n4486,n22,n4485);
not gate_4467(n4487,n4486);
and gate_4468(n4488,n39,n1665);
not gate_4469(n4489,n4488);
and gate_4470(n4490,pi9,n1808);
and gate_4471(n4491,n328,n4490);
not gate_4472(n4492,n4491);
and gate_4473(n4493,n4489,n4492);
not gate_4474(n4494,n4493);
and gate_4475(n4495,pi0,n4494);
not gate_4476(n4496,n4495);
and gate_4477(n4497,n1707,n1731);
and gate_4478(n4498,n2761,n4497);
not gate_4479(n4499,n4498);
and gate_4480(n4500,n4496,n4499);
not gate_4481(n4501,n4500);
and gate_4482(n4502,pi7,n4501);
not gate_4483(n4503,n4502);
and gate_4484(n4504,n709,n715);
not gate_4485(n4505,n4504);
and gate_4486(n4506,n448,n4505);
and gate_4487(n4507,pi0,n4506);
not gate_4488(n4508,n4507);
and gate_4489(n4509,n4503,n4508);
not gate_4490(n4510,n4509);
and gate_4491(n4511,pi2,n4510);
not gate_4492(n4512,n4511);
and gate_4493(n4513,n4487,n4512);
not gate_4494(n4514,n4513);
and gate_4495(n4515,pi5,n4514);
not gate_4496(n4516,n4515);
and gate_4497(n4517,pi0,n3942);
not gate_4498(n4518,n4517);
and gate_4499(n4519,n20,n1759);
not gate_4500(n4520,n4519);
and gate_4501(n4521,n4518,n4520);
not gate_4502(n4522,n4521);
and gate_4503(n4523,n27,n4522);
not gate_4504(n4524,n4523);
and gate_4505(n4525,n2691,n4524);
not gate_4506(n4526,n4525);
and gate_4507(n4527,pi4,n4526);
not gate_4508(n4528,n4527);
and gate_4509(n4529,n27,n2088);
not gate_4510(n4530,n4529);
and gate_4511(n4531,n233,n2775);
not gate_4512(n4532,n4531);
and gate_4513(n4533,n4530,n4532);
and gate_4514(n4534,n766,n4533);
not gate_4515(n4535,n4534);
and gate_4516(n4536,n4528,n4535);
not gate_4517(n4537,n4536);
and gate_4518(n4538,pi2,n4537);
not gate_4519(n4539,n4538);
and gate_4520(n4540,pi3,n509);
not gate_4521(n4541,n4540);
and gate_4522(n4542,n188,n785);
not gate_4523(n4543,n4542);
and gate_4524(n4544,n4541,n4543);
not gate_4525(n4545,n4544);
and gate_4526(n4546,pi8,n4545);
not gate_4527(n4547,n4546);
and gate_4528(n4548,n592,n1732);
not gate_4529(n4549,n4548);
and gate_4530(n4550,n4547,n4549);
not gate_4531(n4551,n4550);
and gate_4532(n4552,pi0,n4551);
not gate_4533(n4553,n4552);
and gate_4534(n4554,n2276,n3309);
not gate_4535(n4555,n4554);
and gate_4536(n4556,n4553,n4555);
not gate_4537(n4557,n4556);
and gate_4538(n4558,n22,n4557);
not gate_4539(n4559,n4558);
and gate_4540(n4560,n4539,n4559);
not gate_4541(n4561,n4560);
and gate_4542(n4562,n25,n4561);
not gate_4543(n4563,n4562);
and gate_4544(n4564,n4516,n4563);
not gate_4545(n4565,n4564);
and gate_4546(n4566,n21,n4565);
not gate_4547(n4567,n4566);
and gate_4548(n4568,n247,n662);
not gate_4549(n4569,n4568);
and gate_4550(n4570,n1177,n4303);
not gate_4551(n4571,n4570);
and gate_4552(n4572,n4569,n4571);
not gate_4553(n4573,n4572);
and gate_4554(n4574,n24,n4573);
not gate_4555(n4575,n4574);
and gate_4556(n4576,n74,n195);
and gate_4557(n4577,n20,n4576);
not gate_4558(n4578,n4577);
and gate_4559(n4579,n4575,n4578);
not gate_4560(n4580,n4579);
and gate_4561(n4581,pi3,n4580);
not gate_4562(n4582,n4581);
and gate_4563(n4583,pi4,n632);
not gate_4564(n4584,n4583);
and gate_4565(n4585,pi0,pi4);
not gate_4566(n4586,n4585);
and gate_4567(n4587,n773,n4586);
not gate_4568(n4588,n4587);
and gate_4569(n4589,n4584,n4588);
and gate_4570(n4590,n960,n4589);
not gate_4571(n4591,n4590);
and gate_4572(n4592,n4582,n4591);
not gate_4573(n4593,n4592);
and gate_4574(n4594,n27,n4593);
not gate_4575(n4595,n4594);
and gate_4576(n4596,n632,n1708);
and gate_4577(n4597,n1175,n4596);
and gate_4578(n4598,pi0,n4597);
not gate_4579(n4599,n4598);
and gate_4580(n4600,n384,n677);
and gate_4581(n4601,n3905,n4600);
not gate_4582(n4602,n4601);
and gate_4583(n4603,n4599,n4602);
not gate_4584(n4604,n4603);
and gate_4585(n4605,n23,n4604);
not gate_4586(n4606,n4605);
and gate_4587(n4607,n708,n2409);
not gate_4588(n4608,n4607);
and gate_4589(n4609,n4606,n4608);
not gate_4590(n4610,n4609);
and gate_4591(n4611,pi7,n4610);
not gate_4592(n4612,n4611);
and gate_4593(n4613,n4595,n4612);
not gate_4594(n4614,n4613);
and gate_4595(n4615,n25,n4614);
not gate_4596(n4616,n4615);
and gate_4597(n4617,n20,n327);
not gate_4598(n4618,n4617);
and gate_4599(n4619,pi3,n4055);
and gate_4600(n4620,n3906,n4619);
not gate_4601(n4621,n4620);
and gate_4602(n4622,n4618,n4621);
not gate_4603(n4623,n4622);
and gate_4604(n4624,n29,n4623);
not gate_4605(n4625,n4624);
and gate_4606(n4626,n2650,n2774);
not gate_4607(n4627,n4626);
and gate_4608(n4628,n4625,n4627);
not gate_4609(n4629,n4628);
and gate_4610(n4630,pi4,n4629);
not gate_4611(n4631,n4630);
and gate_4612(n4632,n182,n729);
and gate_4613(n4633,n1686,n4632);
and gate_4614(n4634,pi0,n4633);
not gate_4615(n4635,n4634);
and gate_4616(n4636,n4631,n4635);
not gate_4617(n4637,n4636);
and gate_4618(n4638,pi2,n4637);
not gate_4619(n4639,n4638);
and gate_4620(n4640,n32,n2552);
and gate_4621(n4641,n2463,n4640);
not gate_4622(n4642,n4641);
and gate_4623(n4643,n4639,n4642);
not gate_4624(n4644,n4643);
and gate_4625(n4645,pi5,n4644);
not gate_4626(n4646,n4645);
and gate_4627(n4647,n4616,n4646);
not gate_4628(n4648,n4647);
and gate_4629(n4649,pi1,n4648);
not gate_4630(n4650,n4649);
and gate_4631(n4651,n4567,n4650);
and gate_4632(n4652,n4474,n4651);
not gate_4633(n4653,n4652);
and gate_4634(n4654,pi6,n4653);
not gate_4635(n4655,n4654);
and gate_4636(n4656,n4453,n4655);
and gate_4637(n4657,n4234,n4656);
not gate_4638(po8,n4657);
and gate_4639(n4659,pi2,n2835);
not gate_4640(n4660,n4659);
and gate_4641(n4661,n131,n2182);
not gate_4642(n4662,n4661);
and gate_4643(n4663,n4660,n4662);
not gate_4644(n4664,n4663);
and gate_4645(n4665,pi9,n4664);
not gate_4646(n4666,n4665);
and gate_4647(n4667,n101,n2276);
not gate_4648(n4668,n4667);
and gate_4649(n4669,n4666,n4668);
not gate_4650(n4670,n4669);
and gate_4651(n4671,pi1,n4670);
not gate_4652(n4672,n4671);
and gate_4653(n4673,n21,n463);
and gate_4654(n4674,n1951,n4673);
not gate_4655(n4675,n4674);
and gate_4656(n4676,n4672,n4675);
not gate_4657(n4677,n4676);
and gate_4658(n4678,n23,n4677);
not gate_4659(n4679,n4678);
and gate_4660(n4680,n27,n39);
and gate_4661(n4681,n3378,n4680);
not gate_4662(n4682,n4681);
and gate_4663(n4683,n360,n1741);
not gate_4664(n4684,n4683);
and gate_4665(n4685,n4682,n4684);
not gate_4666(n4686,n4685);
and gate_4667(n4687,n3006,n4686);
not gate_4668(n4688,n4687);
and gate_4669(n4689,n4679,n4688);
not gate_4670(n4690,n4689);
and gate_4671(n4691,pi0,n4690);
not gate_4672(n4692,n4691);
and gate_4673(n4693,n30,n47);
and gate_4674(n4694,n2629,n4693);
not gate_4675(n4695,n4694);
and gate_4676(n4696,n4692,n4695);
and gate_4677(n4697,n847,n2331);
not gate_4678(n4698,n4697);
and gate_4679(n4699,n20,n945);
and gate_4680(n4700,n1787,n4699);
not gate_4681(n4701,n4700);
and gate_4682(n4702,n1671,n1677);
not gate_4683(n4703,n4702);
and gate_4684(n4704,n995,n4703);
and gate_4685(n4705,n84,n4704);
not gate_4686(n4706,n4705);
and gate_4687(n4707,n4701,n4706);
not gate_4688(n4708,n4707);
and gate_4689(n4709,n4698,n4708);
not gate_4690(n4710,n4709);
and gate_4691(n4711,n26,n582);
and gate_4692(n4712,n568,n4711);
and gate_4693(n4713,pi2,n4712);
not gate_4694(n4714,n4713);
and gate_4695(n4715,pi6,n565);
not gate_4696(n4716,n4715);
and gate_4697(n4717,n2243,n4716);
not gate_4698(n4718,n4717);
and gate_4699(n4719,n22,n4718);
not gate_4700(n4720,n4719);
and gate_4701(n4721,n4714,n4720);
not gate_4702(n4722,n4721);
and gate_4703(n4723,n23,n4722);
not gate_4704(n4724,n4723);
and gate_4705(n4725,n1965,n2225);
not gate_4706(n4726,n4725);
and gate_4707(n4727,n21,n4726);
not gate_4708(n4728,n4727);
and gate_4709(n4729,n32,n1419);
not gate_4710(n4730,n4729);
and gate_4711(n4731,n4728,n4730);
not gate_4712(n4732,n4731);
and gate_4713(n4733,n288,n4732);
not gate_4714(n4734,n4733);
and gate_4715(n4735,n4724,n4734);
not gate_4716(n4736,n4735);
and gate_4717(n4737,n20,n4736);
not gate_4718(n4738,n4737);
and gate_4719(n4739,n634,n1739);
not gate_4720(n4740,n4739);
and gate_4721(n4741,n773,n1214);
not gate_4722(n4742,n4741);
and gate_4723(n4743,n4740,n4742);
not gate_4724(n4744,n4743);
and gate_4725(n4745,n23,n4744);
not gate_4726(n4746,n4745);
and gate_4727(n4747,n30,n565);
not gate_4728(n4748,n4747);
and gate_4729(n4749,n4746,n4748);
not gate_4730(n4750,n4749);
and gate_4731(n4751,n29,n4750);
not gate_4732(n4752,n4751);
and gate_4733(n4753,n26,n1759);
and gate_4734(n4754,n104,n4753);
not gate_4735(n4755,n4754);
and gate_4736(n4756,n4752,n4755);
not gate_4737(n4757,n4756);
and gate_4738(n4758,pi0,n4757);
not gate_4739(n4759,n4758);
and gate_4740(n4760,n4738,n4759);
not gate_4741(n4761,n4760);
and gate_4742(n4762,pi4,n4761);
not gate_4743(n4763,n4762);
and gate_4744(n4764,pi3,n195);
not gate_4745(n4765,n4764);
and gate_4746(n4766,n1911,n4764);
and gate_4747(n4767,pi2,n4766);
not gate_4748(n4768,n4767);
and gate_4749(n4769,n37,n586);
not gate_4750(n4770,n4769);
and gate_4751(n4771,n4768,n4770);
not gate_4752(n4772,n4771);
and gate_4753(n4773,n26,n4772);
not gate_4754(n4774,n4773);
and gate_4755(n4775,n925,n1674);
and gate_4756(n4776,n945,n4775);
not gate_4757(n4777,n4776);
and gate_4758(n4778,n4774,n4777);
not gate_4759(n4779,n4778);
and gate_4760(n4780,pi0,n4779);
not gate_4761(n4781,n4780);
and gate_4762(n4782,n23,n1668);
not gate_4763(n4783,n4782);
and gate_4764(n4784,n1505,n4783);
not gate_4765(n4785,n4784);
and gate_4766(n4786,n29,n4785);
not gate_4767(n4787,n4786);
and gate_4768(n4788,n32,n1506);
not gate_4769(n4789,n4788);
and gate_4770(n4790,n4787,n4789);
not gate_4771(n4791,n4790);
and gate_4772(n4792,pi2,n4791);
not gate_4773(n4793,n4792);
and gate_4774(n4794,pi6,n247);
and gate_4775(n4795,n37,n4794);
not gate_4776(n4796,n4795);
and gate_4777(n4797,n4793,n4796);
not gate_4778(n4798,n4797);
and gate_4779(n4799,n21,n4798);
not gate_4780(n4800,n4799);
and gate_4781(n4801,n247,n874);
not gate_4782(n4802,n4801);
and gate_4783(n4803,n1419,n4801);
not gate_4784(n4804,n4803);
and gate_4785(n4805,n4800,n4804);
not gate_4786(n4806,n4805);
and gate_4787(n4807,n20,n4806);
not gate_4788(n4808,n4807);
and gate_4789(n4809,n4781,n4808);
not gate_4790(n4810,n4809);
and gate_4791(n4811,n24,n4810);
not gate_4792(n4812,n4811);
and gate_4793(n4813,n4763,n4812);
not gate_4794(n4814,n4813);
and gate_4795(n4815,n27,n4814);
not gate_4796(n4816,n4815);
and gate_4797(n4817,n23,n1513);
not gate_4798(n4818,n4817);
and gate_4799(n4819,pi0,n288);
not gate_4800(n4820,n4819);
and gate_4801(n4821,n4818,n4820);
not gate_4802(n4822,n4821);
and gate_4803(n4823,n24,n4822);
not gate_4804(n4824,n4823);
and gate_4805(n4825,n365,n1152);
and gate_4806(n4826,pi0,n4825);
not gate_4807(n4827,n4826);
and gate_4808(n4828,n4824,n4827);
not gate_4809(n4829,n4828);
and gate_4810(n4830,pi1,n4829);
not gate_4811(n4831,n4830);
and gate_4812(n4832,n1649,n3358);
not gate_4813(n4833,n4832);
and gate_4814(n4834,pi6,n4833);
not gate_4815(n4835,n4834);
and gate_4816(n4836,n37,n1154);
not gate_4817(n4837,n4836);
and gate_4818(n4838,n4835,n4837);
not gate_4819(n4839,n4838);
and gate_4820(n4840,n20,n4839);
not gate_4821(n4841,n4840);
and gate_4822(n4842,n712,n3032);
not gate_4823(n4843,n4842);
and gate_4824(n4844,n4841,n4843);
not gate_4825(n4845,n4844);
and gate_4826(n4846,n21,n4845);
not gate_4827(n4847,n4846);
and gate_4828(n4848,n4831,n4847);
not gate_4829(n4849,n4848);
and gate_4830(n4850,pi9,n4849);
not gate_4831(n4851,n4850);
and gate_4832(n4852,n364,n1201);
and gate_4833(n4853,n691,n4852);
and gate_4834(n4854,n24,n4853);
not gate_4835(n4855,n4854);
and gate_4836(n4856,n23,n78);
not gate_4837(n4857,n4856);
and gate_4838(n4858,n4855,n4857);
not gate_4839(n4859,n4858);
and gate_4840(n4860,pi6,n4859);
not gate_4841(n4861,n4860);
and gate_4842(n4862,n106,n644);
and gate_4843(n4863,n531,n4862);
not gate_4844(n4864,n4863);
and gate_4845(n4865,n4861,n4864);
not gate_4846(n4866,n4865);
and gate_4847(n4867,n29,n4866);
not gate_4848(n4868,n4867);
and gate_4849(n4869,n4851,n4868);
not gate_4850(n4870,n4869);
and gate_4851(n4871,pi8,n4870);
not gate_4852(n4872,n4871);
and gate_4853(n4873,n26,n385);
not gate_4854(n4874,n4873);
and gate_4855(n4875,n1071,n4873);
and gate_4856(n4876,n21,n4875);
not gate_4857(n4877,n4876);
and gate_4858(n4878,n945,n1123);
not gate_4859(n4879,n4878);
and gate_4860(n4880,pi4,n4878);
not gate_4861(n4881,n4880);
and gate_4862(n4882,n4877,n4881);
not gate_4863(n4883,n4882);
and gate_4864(n4884,pi0,n4883);
not gate_4865(n4885,n4884);
and gate_4866(n4886,n98,n1123);
not gate_4867(n4887,n4886);
and gate_4868(n4888,n4874,n4887);
not gate_4869(n4889,n4888);
and gate_4870(n4890,n531,n4889);
not gate_4871(n4891,n4890);
and gate_4872(n4892,n4885,n4891);
not gate_4873(n4893,n4892);
and gate_4874(n4894,n22,n4893);
not gate_4875(n4895,n4894);
and gate_4876(n4896,pi0,n578);
not gate_4877(n4897,n4896);
and gate_4878(n4898,n521,n4897);
not gate_4879(n4899,n4898);
and gate_4880(n4900,n1154,n4899);
and gate_4881(n4901,n30,n4900);
not gate_4882(n4902,n4901);
and gate_4883(n4903,n4895,n4902);
not gate_4884(n4904,n4903);
and gate_4885(n4905,n28,n4904);
not gate_4886(n4906,n4905);
and gate_4887(n4907,n4872,n4906);
not gate_4888(n4908,n4907);
and gate_4889(n4909,pi7,n4908);
not gate_4890(n4910,n4909);
and gate_4891(n4911,n4816,n4910);
not gate_4892(n4912,n4911);
and gate_4893(n4913,pi5,n4912);
not gate_4894(n4914,n4913);
and gate_4895(n4915,n37,n762);
not gate_4896(n4916,n4915);
and gate_4897(n4917,n30,n766);
not gate_4898(n4918,n4917);
and gate_4899(n4919,n4916,n4918);
and gate_4900(n4920,n22,n39);
not gate_4901(n4921,n4920);
and gate_4902(n4922,n613,n4921);
not gate_4903(n4923,n4922);
and gate_4904(n4924,n785,n4923);
not gate_4905(n4925,n4924);
and gate_4906(n4926,n4919,n4925);
not gate_4907(n4927,n4926);
and gate_4908(n4928,n26,n4927);
not gate_4909(n4929,n4928);
and gate_4910(n4930,n714,n874);
not gate_4911(n4931,n4930);
and gate_4912(n4932,pi3,n1690);
not gate_4913(n4933,n4932);
and gate_4914(n4934,n23,n1709);
not gate_4915(n4935,n4934);
and gate_4916(n4936,n4933,n4935);
not gate_4917(n4937,n4936);
and gate_4918(n4938,n1174,n4937);
not gate_4919(n4939,n4938);
and gate_4920(n4940,n4931,n4939);
not gate_4921(n4941,n4940);
and gate_4922(n4942,pi6,n4941);
not gate_4923(n4943,n4942);
and gate_4924(n4944,n4929,n4943);
not gate_4925(n4945,n4944);
and gate_4926(n4946,n21,n4945);
not gate_4927(n4947,n4946);
and gate_4928(n4948,n281,n4765);
not gate_4929(n4949,n4948);
and gate_4930(n4950,pi6,n4949);
not gate_4931(n4951,n4950);
and gate_4932(n4952,n39,n1506);
not gate_4933(n4953,n4952);
and gate_4934(n4954,n4951,n4953);
not gate_4935(n4955,n4954);
and gate_4936(n4956,pi2,n4955);
not gate_4937(n4957,n4956);
and gate_4938(n4958,n37,n2515);
not gate_4939(n4959,n4958);
and gate_4940(n4960,n4957,n4959);
not gate_4941(n4961,n4960);
and gate_4942(n4962,n1003,n4961);
not gate_4943(n4963,n4962);
and gate_4944(n4964,n4947,n4963);
not gate_4945(n4965,n4964);
and gate_4946(n4966,pi7,n4965);
not gate_4947(n4967,n4966);
and gate_4948(n4968,n1245,n3137);
not gate_4949(n4969,n4968);
and gate_4950(n4970,n946,n4969);
and gate_4951(n4971,pi2,n4970);
not gate_4952(n4972,n4971);
and gate_4953(n4973,n644,n3139);
not gate_4954(n4974,n4973);
and gate_4955(n4975,n4972,n4974);
not gate_4956(n4976,n4975);
and gate_4957(n4977,n28,n4976);
not gate_4958(n4978,n4977);
and gate_4959(n4979,n21,n1644);
not gate_4960(n4980,n4979);
and gate_4961(n4981,n4879,n4980);
not gate_4962(n4982,n4981);
and gate_4963(n4983,n630,n4982);
not gate_4964(n4984,n4983);
and gate_4965(n4985,n4978,n4984);
not gate_4966(n4986,n4985);
and gate_4967(n4987,pi4,n4986);
not gate_4968(n4988,n4987);
and gate_4969(n4989,n194,n1127);
and gate_4970(n4990,n1912,n4989);
and gate_4971(n4991,n1648,n4990);
not gate_4972(n4992,n4991);
and gate_4973(n4993,n4988,n4992);
not gate_4974(n4994,n4993);
and gate_4975(n4995,n27,n4994);
not gate_4976(n4996,n4995);
and gate_4977(n4997,n4967,n4996);
not gate_4978(n4998,n4997);
and gate_4979(n4999,n20,n4998);
not gate_4980(n5000,n4999);
and gate_4981(n5001,n962,n1321);
not gate_4982(n5002,n5001);
and gate_4983(n5003,n174,n1325);
not gate_4984(n5004,n5003);
and gate_4985(n5005,n5002,n5004);
and gate_4986(n5006,n22,n5005);
not gate_4987(n5007,n5006);
and gate_4988(n5008,n182,n1294);
not gate_4989(n5009,n5008);
and gate_4990(n5010,n874,n5009);
not gate_4991(n5011,n5010);
and gate_4992(n5012,n5007,n5011);
not gate_4993(n5013,n5012);
and gate_4994(n5014,n28,n5013);
not gate_4995(n5015,n5014);
and gate_4996(n5016,n1492,n1587);
not gate_4997(n5017,n5016);
and gate_4998(n5018,n1505,n5017);
and gate_4999(n5019,n636,n5018);
not gate_5000(n5020,n5019);
and gate_5001(n5021,n5015,n5020);
not gate_5002(n5022,n5021);
and gate_5003(n5023,pi1,n5022);
not gate_5004(n5024,n5023);
and gate_5005(n5025,n22,n778);
not gate_5006(n5026,n5025);
and gate_5007(n5027,n4802,n5026);
not gate_5008(n5028,n5027);
and gate_5009(n5029,n1428,n5028);
not gate_5010(n5030,n5029);
and gate_5011(n5031,n5024,n5030);
not gate_5012(n5032,n5031);
and gate_5013(n5033,pi4,n5032);
not gate_5014(n5034,n5033);
and gate_5015(n5035,n30,n3239);
not gate_5016(n5036,n5035);
and gate_5017(n5037,n1200,n3142);
and gate_5018(n5038,n672,n5037);
not gate_5019(n5039,n5038);
and gate_5020(n5040,n5036,n5039);
not gate_5021(n5041,n5040);
and gate_5022(n5042,n28,n5041);
not gate_5023(n5043,n5042);
and gate_5024(n5044,n23,n4681);
not gate_5025(n5045,n5044);
and gate_5026(n5046,n5043,n5045);
not gate_5027(n5047,n5046);
and gate_5028(n5048,pi1,n5047);
not gate_5029(n5049,n5048);
and gate_5030(n5050,n21,n37);
and gate_5031(n5051,n4164,n5050);
not gate_5032(n5052,n5051);
and gate_5033(n5053,n5049,n5052);
not gate_5034(n5054,n5053);
and gate_5035(n5055,n24,n5054);
not gate_5036(n5056,n5055);
and gate_5037(n5057,n5034,n5056);
not gate_5038(n5058,n5057);
and gate_5039(n5059,pi0,n5058);
not gate_5040(n5060,n5059);
and gate_5041(n5061,n5000,n5060);
and gate_5042(n5062,n74,n1964);
not gate_5043(n5063,n5062);
and gate_5044(n5064,n80,n1741);
not gate_5045(n5065,n5064);
and gate_5046(n5066,n5063,n5065);
not gate_5047(n5067,n5066);
and gate_5048(n5068,pi0,n5067);
not gate_5049(n5069,n5068);
and gate_5050(n5070,n20,n165);
and gate_5051(n5071,n41,n5070);
not gate_5052(n5072,n5071);
and gate_5053(n5073,n5069,n5072);
not gate_5054(n5074,n5073);
and gate_5055(n5075,n1483,n5074);
and gate_5056(n5076,n730,n5075);
not gate_5057(n5077,n5076);
and gate_5058(n5078,n5061,n5077);
not gate_5059(n5079,n5078);
and gate_5060(n5080,n25,n5079);
not gate_5061(n5081,n5080);
and gate_5062(n5082,n4914,n5081);
and gate_5063(n5083,n4710,n5082);
and gate_5064(n5084,n4696,n5083);
not gate_5065(po9,n5084);
endmodule
