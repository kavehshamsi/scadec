// Verilog File 
module apex4 (vdd,pi0,pi1,pi2,pi3,pi4,pi5,pi6,pi7,
pi8,po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18);

input vdd,pi0,pi1,pi2,pi3,pi4,pi5,pi6,pi7,
pi8;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18;

wire n28,n30,n31,n32,n33,n34,n35,n36,n37,
n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,
n48,n49,n50,n51,n52,n53,n54,n55,n56,n57,
n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,
n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,
n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,
n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,
n98,n99,n100,n101,n102,n103,n104,n105,n106,n107,
n108,n109,n110,n111,n112,n113,n114,n115,n116,n117,
n118,n119,n120,n121,n122,n123,n124,n125,n126,n127,
n128,n129,n130,n131,n132,n133,n134,n135,n136,n137,
n138,n139,n140,n141,n142,n143,n144,n145,n146,n147,
n148,n149,n150,n151,n152,n153,n154,n155,n156,n157,
n158,n159,n160,n161,n162,n163,n164,n165,n166,n167,
n168,n169,n170,n171,n172,n173,n174,n175,n176,n177,
n178,n179,n180,n181,n182,n183,n184,n185,n186,n187,
n188,n189,n190,n191,n192,n193,n194,n195,n196,n197,
n198,n199,n200,n201,n202,n203,n204,n205,n206,n207,
n208,n209,n210,n211,n212,n213,n214,n215,n216,n217,
n218,n219,n220,n221,n222,n223,n224,n225,n226,n227,
n228,n229,n230,n231,n232,n233,n234,n235,n236,n237,
n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,
n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,
n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,
n268,n269,n270,n271,n272,n273,n274,n275,n276,n277,
n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,
n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,
n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,
n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,
n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,
n329,n330,n331,n332,n333,n334,n335,n336,n337,n338,
n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,
n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,
n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,
n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,
n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,
n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,
n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,
n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,
n419,n420,n421,n422,n423,n424,n425,n426,n427,n428,
n429,n430,n431,n432,n433,n434,n435,n436,n437,n438,
n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,
n449,n450,n451,n452,n453,n454,n455,n456,n457,n458,
n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,
n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,
n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,
n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,
n499,n500,n501,n502,n503,n504,n505,n506,n507,n508,
n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,
n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,
n529,n530,n531,n532,n533,n534,n535,n536,n537,n538,
n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,
n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,
n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,
n569,n570,n571,n572,n573,n574,n575,n576,n577,n578,
n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,
n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,
n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,
n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,
n619,n620,n621,n622,n623,n624,n625,n626,n627,n628,
n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,
n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,
n649,n650,n651,n652,n653,n654,n655,n656,n657,n658,
n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,
n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,
n679,n680,n681,n682,n683,n684,n685,n686,n687,n688,
n689,n690,n691,n692,n693,n694,n695,n696,n697,n698,
n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,
n709,n710,n711,n712,n713,n714,n715,n716,n717,n718,
n719,n720,n721,n722,n723,n724,n725,n726,n727,n728,
n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,
n739,n740,n741,n742,n743,n744,n745,n746,n747,n748,
n749,n750,n751,n752,n753,n754,n755,n756,n757,n758,
n759,n760,n761,n762,n763,n764,n765,n766,n767,n768,
n769,n770,n771,n772,n773,n774,n775,n776,n777,n778,
n779,n780,n781,n782,n783,n784,n785,n786,n787,n788,
n789,n790,n791,n792,n793,n794,n795,n796,n797,n798,
n799,n800,n801,n802,n803,n804,n805,n806,n807,n808,
n809,n811,n812,n813,n814,n815,n816,n817,n818,n819,
n820,n821,n822,n823,n824,n825,n826,n827,n828,n829,
n830,n831,n832,n833,n834,n835,n836,n837,n838,n839,
n840,n841,n842,n843,n844,n845,n846,n847,n848,n849,
n850,n851,n852,n853,n854,n855,n856,n857,n858,n859,
n860,n861,n862,n863,n864,n865,n866,n867,n868,n869,
n870,n871,n872,n873,n874,n875,n876,n877,n878,n879,
n880,n881,n882,n883,n884,n885,n886,n887,n888,n889,
n890,n891,n892,n893,n894,n895,n896,n897,n898,n899,
n900,n901,n902,n903,n904,n905,n906,n907,n908,n909,
n910,n911,n912,n913,n914,n915,n916,n917,n918,n919,
n920,n921,n922,n923,n924,n925,n926,n927,n928,n929,
n930,n931,n932,n933,n934,n935,n936,n937,n938,n939,
n940,n941,n942,n943,n944,n945,n946,n947,n948,n949,
n950,n951,n952,n953,n954,n955,n956,n957,n958,n959,
n960,n961,n962,n963,n964,n965,n966,n967,n968,n969,
n970,n971,n972,n973,n974,n975,n976,n977,n978,n979,
n980,n981,n982,n983,n984,n985,n986,n987,n988,n989,
n990,n991,n992,n993,n994,n995,n996,n997,n998,n999,
n1000,n1001,n1002,n1003,n1004,n1005,n1006,n1007,n1008,n1009,
n1010,n1011,n1012,n1013,n1014,n1015,n1016,n1017,n1018,n1019,
n1020,n1021,n1022,n1023,n1024,n1025,n1026,n1027,n1028,n1029,
n1030,n1031,n1032,n1033,n1034,n1035,n1036,n1037,n1038,n1039,
n1040,n1041,n1042,n1043,n1044,n1045,n1046,n1047,n1048,n1049,
n1050,n1051,n1052,n1053,n1054,n1055,n1056,n1057,n1058,n1059,
n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,n1069,
n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,n1079,
n1080,n1081,n1082,n1083,n1084,n1085,n1086,n1087,n1088,n1089,
n1090,n1091,n1092,n1093,n1094,n1095,n1096,n1097,n1098,n1099,
n1100,n1101,n1102,n1103,n1104,n1105,n1106,n1107,n1108,n1109,
n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,n1118,n1119,
n1120,n1121,n1122,n1123,n1124,n1125,n1126,n1127,n1128,n1129,
n1130,n1131,n1132,n1133,n1134,n1135,n1136,n1137,n1138,n1139,
n1140,n1141,n1142,n1143,n1144,n1145,n1146,n1147,n1148,n1149,
n1150,n1151,n1152,n1153,n1154,n1155,n1156,n1157,n1158,n1159,
n1160,n1161,n1162,n1163,n1164,n1165,n1166,n1167,n1168,n1169,
n1170,n1171,n1172,n1173,n1174,n1175,n1176,n1177,n1178,n1179,
n1180,n1181,n1182,n1183,n1184,n1185,n1186,n1187,n1188,n1189,
n1190,n1191,n1192,n1193,n1194,n1195,n1196,n1197,n1198,n1199,
n1200,n1201,n1202,n1203,n1204,n1205,n1206,n1207,n1208,n1209,
n1210,n1211,n1212,n1213,n1215,n1216,n1217,n1218,n1219,n1220,
n1221,n1222,n1223,n1224,n1225,n1226,n1227,n1228,n1229,n1230,
n1231,n1232,n1233,n1234,n1235,n1236,n1237,n1238,n1239,n1240,
n1241,n1242,n1243,n1244,n1245,n1246,n1247,n1248,n1249,n1250,
n1251,n1252,n1253,n1254,n1255,n1256,n1257,n1258,n1259,n1260,
n1261,n1262,n1263,n1264,n1265,n1266,n1267,n1268,n1269,n1270,
n1271,n1272,n1273,n1274,n1275,n1276,n1277,n1278,n1279,n1280,
n1281,n1282,n1283,n1284,n1285,n1286,n1287,n1288,n1289,n1290,
n1291,n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,n1300,
n1301,n1302,n1303,n1304,n1305,n1306,n1307,n1308,n1309,n1310,
n1311,n1312,n1313,n1314,n1315,n1316,n1317,n1318,n1319,n1320,
n1321,n1322,n1323,n1324,n1325,n1326,n1327,n1328,n1329,n1330,
n1331,n1332,n1333,n1334,n1335,n1336,n1337,n1338,n1339,n1340,
n1341,n1342,n1343,n1344,n1345,n1346,n1347,n1348,n1349,n1350,
n1351,n1352,n1353,n1354,n1355,n1356,n1357,n1358,n1359,n1360,
n1361,n1362,n1363,n1364,n1365,n1366,n1367,n1368,n1369,n1370,
n1371,n1372,n1373,n1374,n1375,n1376,n1377,n1378,n1379,n1380,
n1381,n1382,n1383,n1384,n1385,n1386,n1387,n1388,n1389,n1390,
n1391,n1392,n1393,n1394,n1395,n1396,n1397,n1398,n1399,n1400,
n1401,n1402,n1403,n1404,n1405,n1406,n1407,n1408,n1409,n1410,
n1411,n1412,n1413,n1414,n1415,n1416,n1417,n1418,n1419,n1420,
n1421,n1422,n1423,n1424,n1425,n1426,n1427,n1428,n1429,n1430,
n1431,n1432,n1433,n1434,n1435,n1436,n1437,n1438,n1439,n1440,
n1441,n1442,n1443,n1444,n1445,n1446,n1447,n1448,n1449,n1450,
n1451,n1452,n1453,n1454,n1455,n1456,n1457,n1458,n1459,n1460,
n1461,n1462,n1463,n1464,n1465,n1466,n1467,n1468,n1469,n1470,
n1471,n1472,n1473,n1474,n1475,n1476,n1477,n1478,n1479,n1480,
n1481,n1482,n1483,n1484,n1485,n1486,n1487,n1488,n1489,n1490,
n1491,n1492,n1493,n1494,n1495,n1496,n1497,n1498,n1499,n1500,
n1501,n1502,n1503,n1504,n1505,n1506,n1507,n1508,n1509,n1510,
n1511,n1512,n1513,n1514,n1515,n1516,n1517,n1518,n1519,n1520,
n1521,n1522,n1523,n1524,n1525,n1526,n1527,n1528,n1529,n1530,
n1531,n1532,n1533,n1534,n1535,n1536,n1537,n1538,n1539,n1540,
n1541,n1542,n1543,n1544,n1545,n1546,n1547,n1548,n1549,n1550,
n1551,n1552,n1553,n1554,n1555,n1556,n1557,n1558,n1559,n1560,
n1561,n1562,n1563,n1564,n1565,n1566,n1567,n1568,n1569,n1570,
n1571,n1572,n1573,n1574,n1575,n1576,n1577,n1578,n1579,n1580,
n1581,n1582,n1583,n1584,n1585,n1586,n1587,n1588,n1589,n1590,
n1591,n1592,n1593,n1594,n1595,n1596,n1597,n1598,n1599,n1600,
n1601,n1602,n1603,n1604,n1605,n1606,n1607,n1608,n1609,n1610,
n1611,n1612,n1613,n1614,n1615,n1616,n1617,n1618,n1619,n1620,
n1621,n1622,n1623,n1624,n1625,n1626,n1627,n1628,n1629,n1630,
n1631,n1632,n1633,n1634,n1635,n1636,n1637,n1638,n1639,n1640,
n1641,n1642,n1643,n1644,n1645,n1646,n1647,n1648,n1649,n1650,
n1651,n1652,n1653,n1654,n1655,n1656,n1657,n1658,n1659,n1660,
n1661,n1662,n1663,n1665,n1666,n1667,n1668,n1669,n1670,n1671,
n1672,n1673,n1674,n1675,n1676,n1677,n1678,n1679,n1680,n1681,
n1682,n1683,n1684,n1685,n1686,n1687,n1688,n1689,n1690,n1691,
n1692,n1693,n1694,n1695,n1696,n1697,n1698,n1699,n1700,n1701,
n1702,n1703,n1704,n1705,n1706,n1707,n1708,n1709,n1710,n1711,
n1712,n1713,n1714,n1715,n1716,n1717,n1718,n1719,n1720,n1721,
n1722,n1723,n1724,n1725,n1726,n1727,n1728,n1729,n1730,n1731,
n1732,n1733,n1734,n1735,n1736,n1737,n1738,n1739,n1740,n1741,
n1742,n1743,n1744,n1745,n1746,n1747,n1748,n1749,n1750,n1751,
n1752,n1753,n1754,n1755,n1756,n1757,n1758,n1759,n1760,n1761,
n1762,n1763,n1764,n1765,n1766,n1767,n1768,n1769,n1770,n1771,
n1772,n1773,n1774,n1775,n1776,n1777,n1778,n1779,n1780,n1781,
n1782,n1783,n1784,n1785,n1786,n1787,n1788,n1789,n1790,n1791,
n1792,n1793,n1794,n1795,n1796,n1797,n1798,n1799,n1800,n1801,
n1802,n1803,n1804,n1805,n1806,n1807,n1808,n1809,n1810,n1811,
n1812,n1813,n1814,n1815,n1816,n1817,n1818,n1819,n1820,n1821,
n1822,n1823,n1824,n1825,n1826,n1827,n1828,n1829,n1830,n1831,
n1832,n1833,n1834,n1835,n1836,n1837,n1838,n1839,n1840,n1841,
n1842,n1843,n1844,n1845,n1846,n1847,n1848,n1849,n1850,n1851,
n1852,n1853,n1854,n1855,n1856,n1857,n1858,n1859,n1860,n1861,
n1862,n1863,n1864,n1865,n1866,n1867,n1868,n1869,n1870,n1871,
n1872,n1873,n1874,n1875,n1876,n1877,n1878,n1879,n1880,n1881,
n1882,n1883,n1884,n1885,n1886,n1887,n1888,n1889,n1890,n1891,
n1892,n1893,n1894,n1895,n1896,n1897,n1898,n1899,n1900,n1901,
n1902,n1903,n1904,n1905,n1906,n1907,n1908,n1909,n1910,n1911,
n1912,n1913,n1914,n1915,n1916,n1917,n1918,n1919,n1920,n1921,
n1922,n1923,n1924,n1925,n1926,n1927,n1928,n1929,n1930,n1931,
n1932,n1933,n1934,n1935,n1936,n1937,n1938,n1939,n1940,n1941,
n1942,n1943,n1944,n1945,n1946,n1947,n1948,n1949,n1950,n1951,
n1952,n1953,n1954,n1955,n1956,n1957,n1958,n1959,n1960,n1961,
n1962,n1963,n1964,n1965,n1966,n1967,n1968,n1969,n1970,n1971,
n1972,n1973,n1974,n1975,n1976,n1977,n1978,n1979,n1980,n1981,
n1982,n1983,n1984,n1985,n1986,n1987,n1988,n1989,n1990,n1991,
n1992,n1993,n1994,n1995,n1996,n1997,n1998,n1999,n2000,n2001,
n2002,n2003,n2004,n2005,n2006,n2007,n2008,n2009,n2010,n2011,
n2012,n2013,n2014,n2015,n2016,n2017,n2018,n2019,n2020,n2021,
n2022,n2023,n2024,n2025,n2026,n2027,n2028,n2029,n2030,n2031,
n2032,n2033,n2034,n2035,n2036,n2037,n2038,n2039,n2040,n2041,
n2042,n2043,n2044,n2045,n2046,n2047,n2048,n2049,n2050,n2051,
n2052,n2053,n2054,n2055,n2056,n2057,n2058,n2059,n2060,n2061,
n2062,n2063,n2064,n2065,n2066,n2067,n2068,n2069,n2070,n2071,
n2072,n2073,n2074,n2075,n2076,n2077,n2078,n2079,n2080,n2081,
n2082,n2083,n2084,n2085,n2086,n2087,n2088,n2089,n2090,n2091,
n2093,n2094,n2095,n2096,n2097,n2098,n2099,n2100,n2101,n2102,
n2103,n2104,n2105,n2106,n2107,n2108,n2109,n2110,n2111,n2112,
n2113,n2114,n2115,n2116,n2117,n2118,n2119,n2120,n2121,n2122,
n2123,n2124,n2125,n2126,n2127,n2128,n2129,n2130,n2131,n2132,
n2133,n2134,n2135,n2136,n2137,n2138,n2139,n2140,n2141,n2142,
n2143,n2144,n2145,n2146,n2147,n2148,n2149,n2150,n2151,n2152,
n2153,n2154,n2155,n2156,n2157,n2158,n2159,n2160,n2161,n2162,
n2163,n2164,n2165,n2166,n2167,n2168,n2169,n2170,n2171,n2172,
n2173,n2174,n2175,n2176,n2177,n2178,n2179,n2180,n2181,n2182,
n2183,n2184,n2185,n2186,n2187,n2188,n2189,n2190,n2191,n2192,
n2193,n2194,n2195,n2196,n2197,n2198,n2199,n2200,n2201,n2202,
n2203,n2204,n2205,n2206,n2207,n2208,n2209,n2210,n2211,n2212,
n2213,n2214,n2215,n2216,n2217,n2218,n2219,n2220,n2221,n2222,
n2223,n2224,n2225,n2226,n2227,n2228,n2229,n2230,n2231,n2232,
n2233,n2234,n2235,n2236,n2237,n2238,n2239,n2240,n2241,n2242,
n2243,n2244,n2245,n2246,n2247,n2248,n2249,n2250,n2251,n2252,
n2253,n2254,n2255,n2256,n2257,n2258,n2259,n2260,n2261,n2262,
n2263,n2264,n2265,n2266,n2267,n2268,n2269,n2270,n2271,n2272,
n2273,n2274,n2275,n2276,n2277,n2278,n2279,n2280,n2281,n2282,
n2283,n2284,n2285,n2286,n2287,n2288,n2289,n2290,n2291,n2292,
n2293,n2294,n2295,n2296,n2297,n2298,n2299,n2300,n2301,n2302,
n2303,n2304,n2305,n2306,n2307,n2308,n2309,n2310,n2311,n2312,
n2313,n2314,n2315,n2316,n2317,n2318,n2319,n2320,n2321,n2322,
n2323,n2324,n2325,n2326,n2327,n2328,n2329,n2330,n2331,n2332,
n2333,n2334,n2335,n2336,n2337,n2338,n2339,n2340,n2341,n2342,
n2343,n2344,n2345,n2346,n2347,n2348,n2349,n2350,n2351,n2352,
n2353,n2354,n2355,n2356,n2357,n2358,n2359,n2360,n2361,n2362,
n2363,n2364,n2365,n2366,n2367,n2368,n2369,n2370,n2371,n2372,
n2373,n2374,n2375,n2376,n2377,n2378,n2379,n2380,n2381,n2382,
n2383,n2384,n2385,n2386,n2387,n2388,n2389,n2390,n2391,n2392,
n2393,n2394,n2395,n2396,n2397,n2398,n2399,n2400,n2401,n2402,
n2403,n2404,n2405,n2406,n2407,n2408,n2409,n2410,n2411,n2412,
n2413,n2414,n2415,n2416,n2417,n2418,n2419,n2420,n2421,n2422,
n2423,n2424,n2425,n2426,n2427,n2428,n2429,n2430,n2431,n2432,
n2433,n2434,n2435,n2436,n2437,n2438,n2439,n2440,n2441,n2442,
n2443,n2444,n2445,n2446,n2447,n2448,n2449,n2450,n2451,n2452,
n2453,n2454,n2455,n2456,n2457,n2458,n2459,n2460,n2461,n2462,
n2463,n2464,n2465,n2466,n2467,n2468,n2469,n2470,n2471,n2472,
n2473,n2474,n2475,n2476,n2477,n2478,n2479,n2480,n2481,n2482,
n2483,n2484,n2485,n2486,n2487,n2488,n2489,n2490,n2491,n2492,
n2493,n2494,n2495,n2496,n2497,n2498,n2499,n2500,n2501,n2502,
n2503,n2504,n2505,n2506,n2507,n2508,n2509,n2510,n2511,n2512,
n2513,n2514,n2515,n2516,n2517,n2518,n2519,n2520,n2521,n2522,
n2523,n2524,n2525,n2526,n2527,n2528,n2529,n2530,n2531,n2532,
n2533,n2534,n2535,n2536,n2537,n2538,n2539,n2540,n2541,n2542,
n2543,n2544,n2545,n2546,n2547,n2548,n2549,n2550,n2551,n2552,
n2553,n2554,n2555,n2556,n2557,n2558,n2559,n2560,n2561,n2562,
n2563,n2564,n2565,n2566,n2567,n2568,n2569,n2570,n2571,n2572,
n2573,n2574,n2575,n2576,n2577,n2579,n2580,n2581,n2582,n2583,
n2584,n2585,n2586,n2587,n2588,n2589,n2590,n2591,n2592,n2593,
n2594,n2595,n2596,n2597,n2598,n2599,n2600,n2601,n2602,n2603,
n2604,n2605,n2606,n2607,n2608,n2609,n2610,n2611,n2612,n2613,
n2614,n2615,n2616,n2617,n2618,n2619,n2620,n2621,n2622,n2623,
n2624,n2625,n2626,n2627,n2628,n2629,n2630,n2631,n2632,n2633,
n2634,n2635,n2636,n2637,n2638,n2639,n2640,n2641,n2642,n2643,
n2644,n2645,n2646,n2647,n2648,n2649,n2650,n2651,n2652,n2653,
n2654,n2655,n2656,n2657,n2658,n2659,n2660,n2661,n2662,n2663,
n2664,n2665,n2666,n2667,n2668,n2669,n2670,n2671,n2672,n2673,
n2674,n2675,n2676,n2677,n2678,n2679,n2680,n2681,n2682,n2683,
n2684,n2685,n2686,n2687,n2688,n2689,n2690,n2691,n2692,n2693,
n2694,n2695,n2696,n2697,n2698,n2699,n2700,n2701,n2702,n2703,
n2704,n2705,n2706,n2707,n2708,n2709,n2710,n2711,n2712,n2713,
n2714,n2715,n2716,n2717,n2718,n2719,n2720,n2721,n2722,n2723,
n2724,n2725,n2726,n2727,n2728,n2729,n2730,n2731,n2732,n2733,
n2734,n2735,n2736,n2737,n2738,n2739,n2740,n2741,n2742,n2743,
n2744,n2745,n2746,n2747,n2748,n2749,n2750,n2751,n2752,n2753,
n2754,n2755,n2756,n2757,n2758,n2759,n2760,n2761,n2762,n2763,
n2764,n2765,n2766,n2767,n2768,n2769,n2770,n2771,n2772,n2773,
n2774,n2775,n2776,n2777,n2778,n2779,n2780,n2781,n2782,n2783,
n2784,n2785,n2786,n2787,n2788,n2789,n2790,n2791,n2792,n2793,
n2794,n2795,n2796,n2797,n2798,n2799,n2800,n2801,n2802,n2803,
n2804,n2805,n2806,n2807,n2808,n2809,n2810,n2811,n2812,n2813,
n2814,n2815,n2816,n2817,n2818,n2819,n2820,n2821,n2822,n2823,
n2824,n2825,n2826,n2827,n2828,n2829,n2830,n2831,n2832,n2833,
n2834,n2835,n2836,n2837,n2838,n2839,n2840,n2841,n2842,n2843,
n2844,n2845,n2846,n2847,n2848,n2849,n2850,n2851,n2852,n2853,
n2854,n2855,n2856,n2857,n2858,n2859,n2860,n2861,n2862,n2863,
n2864,n2865,n2866,n2867,n2868,n2869,n2870,n2871,n2872,n2873,
n2874,n2875,n2876,n2877,n2878,n2879,n2880,n2881,n2882,n2883,
n2884,n2885,n2886,n2887,n2888,n2889,n2890,n2891,n2892,n2893,
n2894,n2895,n2896,n2897,n2898,n2899,n2900,n2901,n2902,n2903,
n2904,n2905,n2906,n2907,n2908,n2909,n2910,n2911,n2912,n2913,
n2914,n2915,n2916,n2917,n2918,n2919,n2920,n2921,n2922,n2923,
n2924,n2925,n2926,n2927,n2928,n2929,n2930,n2931,n2932,n2933,
n2934,n2935,n2936,n2937,n2938,n2939,n2940,n2941,n2942,n2943,
n2944,n2945,n2946,n2947,n2948,n2949,n2950,n2951,n2952,n2953,
n2954,n2955,n2956,n2957,n2958,n2959,n2960,n2961,n2962,n2963,
n2964,n2965,n2966,n2967,n2968,n2969,n2970,n2971,n2972,n2973,
n2974,n2975,n2976,n2977,n2978,n2979,n2980,n2981,n2982,n2983,
n2984,n2985,n2986,n2987,n2988,n2989,n2990,n2991,n2992,n2993,
n2994,n2995,n2996,n2997,n2998,n2999,n3000,n3001,n3002,n3003,
n3004,n3005,n3006,n3007,n3008,n3009,n3010,n3011,n3012,n3013,
n3014,n3015,n3016,n3017,n3018,n3019,n3021,n3022,n3023,n3024,
n3025,n3026,n3027,n3028,n3029,n3030,n3031,n3032,n3033,n3034,
n3035,n3036,n3037,n3038,n3039,n3040,n3041,n3042,n3043,n3044,
n3045,n3046,n3047,n3048,n3049,n3050,n3051,n3052,n3053,n3054,
n3055,n3056,n3057,n3058,n3059,n3060,n3061,n3062,n3063,n3064,
n3065,n3066,n3067,n3068,n3069,n3070,n3071,n3072,n3073,n3074,
n3075,n3076,n3077,n3078,n3079,n3080,n3081,n3082,n3083,n3084,
n3085,n3086,n3087,n3088,n3089,n3090,n3091,n3092,n3093,n3094,
n3095,n3096,n3097,n3098,n3099,n3100,n3101,n3102,n3103,n3104,
n3105,n3106,n3107,n3108,n3109,n3110,n3111,n3112,n3113,n3114,
n3115,n3116,n3117,n3118,n3119,n3120,n3121,n3122,n3123,n3124,
n3125,n3126,n3127,n3128,n3129,n3130,n3131,n3132,n3133,n3134,
n3135,n3136,n3137,n3138,n3139,n3140,n3141,n3142,n3143,n3144,
n3145,n3146,n3147,n3148,n3149,n3150,n3151,n3152,n3153,n3154,
n3155,n3156,n3157,n3158,n3159,n3160,n3161,n3162,n3163,n3164,
n3165,n3166,n3167,n3168,n3169,n3170,n3171,n3172,n3173,n3174,
n3175,n3176,n3177,n3178,n3179,n3180,n3181,n3182,n3183,n3184,
n3185,n3186,n3187,n3188,n3189,n3190,n3191,n3192,n3193,n3194,
n3195,n3196,n3197,n3198,n3199,n3200,n3201,n3202,n3203,n3204,
n3205,n3206,n3207,n3208,n3209,n3210,n3211,n3212,n3213,n3214,
n3215,n3216,n3217,n3218,n3219,n3220,n3221,n3222,n3223,n3224,
n3225,n3226,n3227,n3228,n3229,n3230,n3231,n3232,n3233,n3234,
n3235,n3236,n3237,n3238,n3239,n3240,n3241,n3242,n3243,n3244,
n3245,n3246,n3247,n3248,n3249,n3250,n3251,n3252,n3253,n3254,
n3255,n3256,n3257,n3258,n3259,n3260,n3261,n3262,n3263,n3264,
n3265,n3266,n3267,n3268,n3269,n3270,n3271,n3272,n3273,n3274,
n3275,n3276,n3277,n3278,n3279,n3280,n3281,n3282,n3283,n3284,
n3285,n3286,n3287,n3288,n3289,n3290,n3291,n3292,n3293,n3294,
n3295,n3296,n3297,n3298,n3299,n3300,n3301,n3302,n3303,n3304,
n3305,n3306,n3307,n3308,n3309,n3310,n3311,n3312,n3313,n3314,
n3315,n3316,n3317,n3318,n3319,n3320,n3321,n3322,n3323,n3324,
n3325,n3326,n3327,n3328,n3329,n3330,n3331,n3332,n3333,n3334,
n3335,n3336,n3337,n3338,n3339,n3340,n3341,n3342,n3343,n3344,
n3345,n3346,n3347,n3348,n3349,n3350,n3351,n3352,n3353,n3354,
n3355,n3356,n3357,n3358,n3359,n3360,n3361,n3362,n3363,n3364,
n3365,n3366,n3367,n3368,n3369,n3370,n3371,n3372,n3373,n3374,
n3375,n3376,n3377,n3378,n3379,n3380,n3381,n3382,n3383,n3384,
n3385,n3386,n3387,n3388,n3389,n3390,n3391,n3392,n3393,n3394,
n3395,n3396,n3397,n3398,n3399,n3400,n3401,n3402,n3403,n3404,
n3405,n3406,n3407,n3408,n3409,n3411,n3412,n3413,n3414,n3415,
n3416,n3417,n3418,n3419,n3420,n3421,n3422,n3423,n3424,n3425,
n3426,n3427,n3428,n3429,n3430,n3431,n3432,n3433,n3434,n3435,
n3436,n3437,n3438,n3439,n3440,n3441,n3442,n3443,n3444,n3445,
n3446,n3447,n3448,n3449,n3450,n3451,n3452,n3453,n3454,n3455,
n3456,n3457,n3458,n3459,n3460,n3461,n3462,n3463,n3464,n3465,
n3466,n3467,n3468,n3469,n3470,n3471,n3472,n3473,n3474,n3475,
n3476,n3477,n3478,n3479,n3480,n3481,n3482,n3483,n3484,n3485,
n3486,n3487,n3488,n3489,n3490,n3491,n3492,n3493,n3494,n3495,
n3496,n3497,n3498,n3499,n3500,n3501,n3502,n3503,n3504,n3505,
n3506,n3507,n3508,n3509,n3510,n3511,n3512,n3513,n3514,n3515,
n3516,n3517,n3518,n3519,n3520,n3521,n3522,n3523,n3524,n3525,
n3526,n3527,n3528,n3529,n3530,n3531,n3532,n3533,n3534,n3535,
n3536,n3537,n3538,n3539,n3540,n3541,n3542,n3543,n3544,n3545,
n3546,n3547,n3548,n3549,n3550,n3551,n3552,n3553,n3554,n3555,
n3556,n3557,n3558,n3559,n3560,n3561,n3562,n3563,n3564,n3565,
n3566,n3567,n3568,n3569,n3570,n3571,n3572,n3573,n3574,n3575,
n3576,n3577,n3578,n3579,n3580,n3581,n3582,n3583,n3584,n3585,
n3586,n3587,n3588,n3589,n3590,n3591,n3592,n3593,n3594,n3595,
n3596,n3597,n3598,n3599,n3600,n3601,n3602,n3603,n3604,n3605,
n3606,n3607,n3608,n3609,n3610,n3611,n3612,n3613,n3614,n3615,
n3616,n3617,n3618,n3619,n3620,n3621,n3622,n3623,n3624,n3625,
n3626,n3627,n3628,n3629,n3630,n3631,n3632,n3633,n3634,n3635,
n3636,n3637,n3638,n3639,n3640,n3641,n3642,n3643,n3644,n3645,
n3646,n3647,n3648,n3649,n3650,n3651,n3652,n3653,n3654,n3655,
n3656,n3657,n3658,n3659,n3660,n3661,n3662,n3663,n3664,n3665,
n3666,n3667,n3668,n3669,n3670,n3671,n3672,n3673,n3674,n3675,
n3676,n3677,n3678,n3679,n3680,n3681,n3682,n3683,n3684,n3685,
n3686,n3687,n3688,n3689,n3690,n3691,n3692,n3693,n3694,n3695,
n3696,n3697,n3698,n3699,n3700,n3701,n3702,n3703,n3704,n3705,
n3706,n3707,n3708,n3709,n3710,n3711,n3712,n3713,n3714,n3715,
n3716,n3717,n3718,n3719,n3720,n3721,n3722,n3723,n3724,n3725,
n3726,n3727,n3728,n3729,n3730,n3731,n3732,n3733,n3734,n3735,
n3736,n3737,n3738,n3739,n3740,n3741,n3742,n3743,n3744,n3745,
n3746,n3747,n3748,n3749,n3750,n3751,n3752,n3753,n3754,n3755,
n3756,n3757,n3758,n3759,n3760,n3761,n3762,n3763,n3764,n3765,
n3766,n3767,n3768,n3769,n3770,n3771,n3772,n3773,n3774,n3775,
n3776,n3777,n3778,n3779,n3780,n3781,n3782,n3783,n3784,n3785,
n3786,n3787,n3788,n3789,n3790,n3791,n3792,n3793,n3794,n3795,
n3796,n3797,n3798,n3799,n3800,n3801,n3802,n3803,n3804,n3805,
n3806,n3807,n3808,n3809,n3810,n3811,n3812,n3813,n3814,n3815,
n3816,n3817,n3818,n3819,n3820,n3821,n3822,n3823,n3824,n3825,
n3826,n3827,n3828,n3830,n3831,n3832,n3833,n3834,n3835,n3836,
n3837,n3838,n3839,n3840,n3841,n3842,n3843,n3844,n3845,n3846,
n3847,n3848,n3849,n3850,n3851,n3852,n3853,n3854,n3855,n3856,
n3857,n3858,n3859,n3860,n3861,n3862,n3863,n3864,n3865,n3866,
n3867,n3868,n3869,n3870,n3871,n3872,n3873,n3874,n3875,n3876,
n3877,n3878,n3879,n3880,n3881,n3882,n3883,n3884,n3885,n3886,
n3887,n3888,n3889,n3890,n3891,n3892,n3893,n3894,n3895,n3896,
n3897,n3898,n3899,n3900,n3901,n3902,n3903,n3904,n3905,n3906,
n3907,n3908,n3909,n3910,n3911,n3912,n3913,n3914,n3915,n3916,
n3917,n3918,n3919,n3920,n3921,n3922,n3923,n3924,n3925,n3926,
n3927,n3928,n3929,n3930,n3931,n3932,n3933,n3934,n3935,n3936,
n3937,n3938,n3939,n3940,n3941,n3942,n3943,n3944,n3945,n3946,
n3947,n3948,n3949,n3950,n3951,n3952,n3953,n3954,n3955,n3956,
n3957,n3958,n3959,n3960,n3961,n3962,n3963,n3964,n3965,n3966,
n3967,n3968,n3969,n3970,n3971,n3972,n3973,n3974,n3975,n3976,
n3977,n3978,n3979,n3980,n3981,n3982,n3983,n3984,n3985,n3986,
n3987,n3988,n3989,n3990,n3991,n3992,n3993,n3994,n3995,n3996,
n3997,n3998,n3999,n4000,n4001,n4002,n4003,n4004,n4005,n4006,
n4007,n4008,n4009,n4010,n4011,n4012,n4013,n4014,n4015,n4016,
n4017,n4018,n4019,n4020,n4021,n4022,n4023,n4024,n4025,n4026,
n4027,n4028,n4029,n4030,n4031,n4032,n4033,n4034,n4035,n4036,
n4037,n4038,n4039,n4040,n4041,n4042,n4043,n4044,n4045,n4046,
n4047,n4048,n4049,n4050,n4051,n4052,n4053,n4054,n4055,n4056,
n4057,n4058,n4059,n4060,n4061,n4062,n4063,n4064,n4065,n4066,
n4067,n4068,n4069,n4070,n4071,n4072,n4073,n4074,n4075,n4076,
n4077,n4078,n4079,n4080,n4081,n4082,n4083,n4084,n4085,n4086,
n4087,n4088,n4089,n4090,n4091,n4092,n4093,n4094,n4095,n4096,
n4097,n4098,n4099,n4100,n4101,n4102,n4103,n4104,n4105,n4106,
n4107,n4108,n4109,n4110,n4111,n4112,n4113,n4114,n4115,n4116,
n4117,n4118,n4119,n4120,n4121,n4122,n4123,n4124,n4125,n4126,
n4127,n4128,n4129,n4130,n4131,n4132,n4133,n4134,n4135,n4136,
n4137,n4138,n4139,n4140,n4141,n4142,n4143,n4144,n4145,n4146,
n4147,n4148,n4149,n4150,n4151,n4152,n4153,n4154,n4155,n4156,
n4157,n4158,n4159,n4160,n4161,n4162,n4163,n4164,n4165,n4166,
n4167,n4168,n4169,n4170,n4171,n4172,n4173,n4174,n4175,n4176,
n4177,n4178,n4179,n4180,n4181,n4182,n4183,n4184,n4185,n4186,
n4187,n4188,n4189,n4190,n4191,n4192,n4193,n4194,n4195,n4196,
n4197,n4199,n4200,n4201,n4202,n4203,n4204,n4205,n4206,n4207,
n4208,n4209,n4210,n4211,n4212,n4213,n4214,n4215,n4216,n4217,
n4218,n4219,n4220,n4221,n4222,n4223,n4224,n4225,n4226,n4227,
n4228,n4229,n4230,n4231,n4232,n4233,n4234,n4235,n4236,n4237,
n4238,n4239,n4240,n4241,n4242,n4243,n4244,n4245,n4246,n4247,
n4248,n4249,n4250,n4251,n4252,n4253,n4254,n4255,n4256,n4257,
n4258,n4259,n4260,n4261,n4262,n4263,n4264,n4265,n4266,n4267,
n4268,n4269,n4270,n4271,n4272,n4273,n4274,n4275,n4276,n4277,
n4278,n4279,n4280,n4281,n4282,n4283,n4284,n4285,n4286,n4287,
n4288,n4289,n4290,n4291,n4292,n4293,n4294,n4295,n4296,n4297,
n4298,n4299,n4300,n4301,n4302,n4303,n4304,n4305,n4306,n4307,
n4308,n4309,n4310,n4311,n4312,n4313,n4314,n4315,n4316,n4317,
n4318,n4319,n4320,n4321,n4322,n4323,n4324,n4325,n4326,n4327,
n4328,n4329,n4330,n4331,n4332,n4333,n4334,n4335,n4336,n4337,
n4338,n4339,n4340,n4341,n4342,n4343,n4344,n4345,n4346,n4347,
n4348,n4349,n4350,n4351,n4352,n4353,n4354,n4355,n4356,n4357,
n4358,n4359,n4360,n4361,n4362,n4363,n4364,n4365,n4366,n4367,
n4368,n4369,n4370,n4371,n4372,n4373,n4374,n4375,n4376,n4377,
n4378,n4379,n4380,n4381,n4382,n4383,n4384,n4385,n4386,n4387,
n4388,n4389,n4390,n4391,n4392,n4393,n4394,n4395,n4396,n4397,
n4398,n4399,n4400,n4401,n4402,n4403,n4404,n4405,n4406,n4407,
n4408,n4409,n4410,n4411,n4412,n4413,n4414,n4415,n4416,n4417,
n4418,n4419,n4420,n4421,n4422,n4423,n4424,n4425,n4426,n4427,
n4428,n4429,n4430,n4431,n4432,n4433,n4434,n4435,n4436,n4437,
n4438,n4439,n4440,n4441,n4442,n4443,n4444,n4445,n4446,n4447,
n4448,n4449,n4450,n4451,n4452,n4453,n4454,n4455,n4456,n4457,
n4458,n4459,n4460,n4461,n4462,n4463,n4464,n4465,n4466,n4467,
n4468,n4469,n4470,n4471,n4472,n4473,n4475,n4476,n4477,n4478,
n4479,n4480,n4481,n4482,n4483,n4484,n4485,n4486,n4487,n4488,
n4489,n4490,n4491,n4492,n4493,n4494,n4495,n4496,n4497,n4498,
n4499,n4500,n4501,n4502,n4503,n4504,n4505,n4506,n4507,n4508,
n4509,n4510,n4511,n4512,n4513,n4514,n4515,n4516,n4517,n4518,
n4519,n4520,n4521,n4522,n4523,n4524,n4525,n4526,n4527,n4528,
n4529,n4530,n4531,n4532,n4533,n4534,n4535,n4536,n4537,n4538,
n4539,n4540,n4541,n4542,n4543,n4544,n4545,n4546,n4547,n4548,
n4549,n4550,n4551,n4552,n4553,n4554,n4555,n4556,n4557,n4558,
n4559,n4560,n4561,n4562,n4563,n4564,n4565,n4566,n4567,n4568,
n4569,n4570,n4571,n4572,n4573,n4574,n4575,n4576,n4577,n4578,
n4579,n4580,n4581,n4582,n4583,n4584,n4585,n4586,n4587,n4588,
n4589,n4590,n4591,n4592,n4593,n4594,n4595,n4596,n4597,n4598,
n4599,n4600,n4601,n4602,n4603,n4604,n4605,n4606,n4607,n4608,
n4609,n4610,n4611,n4612,n4613,n4614,n4615,n4616,n4617,n4618,
n4619,n4620,n4621,n4622,n4623,n4624,n4625,n4626,n4627,n4628,
n4629,n4630,n4631,n4632,n4633,n4634,n4635,n4636,n4637,n4638,
n4639,n4640,n4641,n4642,n4643,n4644,n4645,n4646,n4647,n4648,
n4649,n4650,n4651,n4652,n4653,n4654,n4655,n4656,n4657,n4658,
n4659,n4660,n4661,n4662,n4663,n4664,n4665,n4666,n4667,n4668,
n4669,n4670,n4671,n4672,n4673,n4674,n4675,n4676,n4678,n4679,
n4680,n4681,n4682,n4683,n4684,n4685,n4686,n4687,n4688,n4689,
n4690,n4691,n4692,n4693,n4694,n4695,n4696,n4697,n4698,n4699,
n4700,n4701,n4702,n4703,n4704,n4705,n4706,n4707,n4708,n4709,
n4710,n4711,n4712,n4713,n4714,n4715,n4716,n4717,n4718,n4719,
n4720,n4721,n4722,n4723,n4724,n4725,n4726,n4727,n4728,n4729,
n4730,n4731,n4732,n4733,n4734,n4735,n4736,n4737,n4738,n4739,
n4740,n4741,n4742,n4743,n4744,n4745,n4746,n4747,n4748,n4749,
n4750,n4751,n4752,n4753,n4754,n4755,n4756,n4757,n4758,n4759,
n4760,n4761,n4762,n4763,n4764,n4765,n4766,n4767,n4768,n4769,
n4770,n4771,n4772,n4773,n4774,n4775,n4776,n4777,n4778,n4779,
n4780,n4781,n4782,n4783,n4784,n4785,n4786,n4787,n4788,n4789,
n4790,n4791,n4792,n4793,n4794,n4795,n4796,n4797,n4798,n4799,
n4800,n4801,n4802,n4803,n4804,n4805,n4806,n4807,n4808,n4809,
n4810,n4811,n4812,n4813,n4814,n4815,n4816,n4817,n4818,n4819,
n4820,n4821,n4822,n4823,n4824,n4825,n4826,n4827,n4828,n4829,
n4830,n4831,n4832,n4833,n4834,n4835,n4836,n4837,n4838,n4839,
n4840,n4841,n4842,n4843,n4844,n4845,n4846,n4847,n4848,n4849,
n4850,n4851,n4852,n4853,n4854,n4855,n4856,n4857,n4858,n4859,
n4860,n4861,n4862,n4863,n4864,n4865,n4866,n4867,n4868,n4869,
n4870,n4871,n4872,n4873,n4874,n4875,n4876,n4877,n4878,n4879,
n4881,n4882,n4883,n4884,n4885,n4886,n4887,n4888,n4889,n4890,
n4891,n4892,n4893,n4894,n4895,n4896,n4897,n4898,n4899,n4900,
n4901,n4902,n4903,n4904,n4905,n4906,n4907,n4908,n4909,n4910,
n4911,n4912,n4913,n4914,n4915,n4916,n4917,n4918,n4919,n4920,
n4921,n4922,n4923,n4924,n4925,n4926,n4927,n4928,n4929,n4930,
n4931,n4932,n4933,n4934,n4935,n4936,n4937,n4938,n4939,n4940,
n4941,n4942,n4943,n4944,n4945,n4946,n4947,n4948,n4949,n4950,
n4951,n4952,n4953,n4954,n4955,n4956,n4957,n4958,n4959,n4960,
n4961,n4962,n4963,n4964,n4965,n4966,n4967,n4968,n4969,n4970,
n4971,n4972,n4973,n4974,n4975,n4976,n4977,n4978,n4979,n4980,
n4981,n4982,n4983,n4984,n4985,n4986,n4987,n4988,n4989,n4990,
n4991,n4992,n4993,n4994,n4995,n4996,n4997,n4998,n4999,n5000,
n5001,n5002,n5003,n5004,n5005,n5006,n5007,n5008,n5009,n5010,
n5011,n5012,n5013,n5014,n5015,n5016,n5017,n5018,n5019,n5020,
n5021,n5022,n5023,n5024,n5025,n5026,n5027,n5028,n5029,n5030,
n5031,n5032,n5033,n5034,n5035,n5036,n5037,n5038,n5039,n5040,
n5041,n5042,n5043,n5044,n5045,n5046,n5047,n5048,n5049,n5050,
n5051,n5052,n5053,n5054,n5055,n5056,n5057,n5058,n5059,n5060,
n5061,n5062,n5063,n5064,n5065,n5066,n5067,n5068,n5069,n5070,
n5071,n5072,n5073,n5074,n5075,n5076,n5077,n5078,n5079,n5080,
n5081,n5082,n5083,n5084,n5085,n5086,n5087,n5088,n5089,n5090,
n5091,n5092,n5093,n5094,n5095,n5096,n5097,n5098,n5099,n5100,
n5101,n5102,n5103,n5104,n5105,n5106,n5107,n5108,n5109,n5110,
n5111,n5112,n5113,n5114,n5115,n5116,n5117,n5118,n5119,n5120,
n5121,n5122,n5123,n5124,n5125,n5126,n5127,n5128,n5129,n5130,
n5131,n5132,n5133,n5134,n5135,n5136,n5137,n5138,n5139,n5140,
n5141,n5142,n5143,n5144,n5145,n5146,n5147,n5148,n5149,n5150,
n5152,n5153,n5154,n5155,n5156,n5157,n5158,n5159,n5160,n5161,
n5162,n5163,n5164,n5165,n5166,n5167,n5168,n5169,n5170,n5171,
n5172,n5173,n5174,n5175,n5176,n5177,n5178,n5179,n5180,n5181,
n5182,n5183,n5184,n5185,n5186,n5187,n5188,n5189,n5190,n5191,
n5192,n5193,n5194,n5195,n5196,n5197,n5198,n5199,n5200,n5201,
n5202,n5203,n5204,n5205,n5206,n5207,n5208,n5209,n5210,n5211,
n5212,n5213,n5214,n5215,n5216,n5217,n5218,n5219,n5220,n5221,
n5222,n5223,n5224,n5225,n5227,n5228,n5229,n5230,n5231,n5232,
n5233,n5234,n5235,n5236,n5237,n5238,n5239,n5240,n5241,n5242,
n5243,n5244,n5245,n5246,n5247,n5248,n5249,n5250,n5251,n5252,
n5253,n5254,n5255,n5256,n5257,n5258,n5259,n5260,n5261,n5262,
n5263,n5264,n5265,n5266,n5267,n5268,n5269,n5270,n5271,n5272,
n5273,n5274,n5275,n5276,n5277,n5278,n5279,n5280,n5281,n5282,
n5283,n5284,n5285,n5287,n5288,n5289,n5290,n5291,n5292,n5293,
n5294,n5295,n5296,n5297,n5298,n5299,n5300,n5301,n5302,n5303,
n5304,n5305,n5306,n5307,n5308,n5309,n5310,n5311,n5312,n5313,
n5314,n5315,n5316,n5317,n5318,n5319,n5320,n5321,n5323,n5324,
n5325,n5326,n5327,n5328,n5329,n5330,n5331,n5332,n5333,n5334,
n5335,n5336,n5337,n5338,n5339,n5340,n5341,n5342,n5343,n5344,
n5345,n5346,n5347,n5348,n5349,n5350,n5351,n5352,n5353,n5354,
n5355,n5356,n5357,n5358,n5359,n5360,n5361,n5362,n5363,n5364,
n5365,n5366,n5367,n5368,n5369,n5370,n5371,n5372,n5373,n5374,
n5375,n5376,n5377,n5378,n5379,n5380,n5381,n5382,n5383,n5384,
n5385,n5386;
vdd);
not gate_1(po00,n28);
not gate_2(n30,pi0);
not gate_3(n31,pi1);
not gate_4(n32,pi2);
not gate_5(n33,pi3);
not gate_6(n34,pi4);
not gate_7(n35,pi5);
not gate_8(n36,pi6);
not gate_9(n37,pi7);
not gate_10(n38,pi8);
and gate_11(n39,pi7,pi8);
not gate_12(n40,n39);
and gate_13(n41,n36,n39);
not gate_14(n42,n41);
and gate_15(n43,n37,n38);
not gate_16(n44,n43);
and gate_17(n45,pi6,n43);
not gate_18(n46,n45);
and gate_19(n47,n42,n46);
not gate_20(n48,n47);
and gate_21(n49,pi3,n48);
not gate_22(n50,n49);
and gate_23(n51,n33,pi6);
not gate_24(n52,n51);
and gate_25(n53,pi7,n38);
not gate_26(n54,n53);
and gate_27(n55,n51,n53);
not gate_28(n56,n55);
and gate_29(n57,n50,n56);
not gate_30(n58,n57);
and gate_31(n59,n30,n58);
not gate_32(n60,n59);
and gate_33(n61,pi7,n54);
not gate_34(n62,n61);
and gate_35(n63,pi6,n62);
not gate_36(n64,n63);
and gate_37(n65,n36,n43);
not gate_38(n66,n65);
and gate_39(n67,n64,n66);
not gate_40(n68,n67);
and gate_41(n69,pi0,n33);
not gate_42(n70,n69);
and gate_43(n71,n68,n69);
not gate_44(n72,n71);
and gate_45(n73,n60,n72);
not gate_46(n74,n73);
and gate_47(n75,pi5,n74);
not gate_48(n76,n75);
and gate_49(n77,pi7,n40);
not gate_50(n78,n77);
and gate_51(n79,pi0,n78);
not gate_52(n80,n79);
and gate_53(n81,n37,pi8);
not gate_54(n82,n81);
and gate_55(n83,n30,n81);
not gate_56(n84,n83);
and gate_57(n85,n80,n84);
not gate_58(n86,n85);
and gate_59(n87,n35,pi6);
not gate_60(n88,n87);
and gate_61(n89,n33,n87);
not gate_62(n90,n89);
and gate_63(n91,n86,n89);
not gate_64(n92,n91);
and gate_65(n93,n76,n92);
not gate_66(n94,n93);
and gate_67(n95,n34,n94);
not gate_68(n96,n95);
and gate_69(n97,n36,n37);
not gate_70(n98,n97);
and gate_71(n99,n35,pi8);
not gate_72(n100,n99);
and gate_73(n101,n97,n100);
and gate_74(n102,pi0,n101);
not gate_75(n103,n102);
and gate_76(n104,pi6,pi7);
not gate_77(n105,n104);
and gate_78(n106,n35,n104);
not gate_79(n107,n106);
and gate_80(n108,n30,n106);
not gate_81(n109,n108);
and gate_82(n110,n103,n109);
not gate_83(n111,n110);
and gate_84(n112,n33,n111);
not gate_85(n113,n112);
and gate_86(n114,pi3,pi5);
not gate_87(n115,n114);
and gate_88(n116,n30,n114);
and gate_89(n117,pi6,n53);
not gate_90(n118,n117);
and gate_91(n119,n116,n117);
not gate_92(n120,n119);
and gate_93(n121,n113,n120);
not gate_94(n122,n121);
and gate_95(n123,pi4,n122);
not gate_96(n124,n123);
and gate_97(n125,n96,n124);
not gate_98(n126,n125);
and gate_99(n127,pi2,n126);
not gate_100(n128,n127);
and gate_101(n129,n35,n81);
not gate_102(n130,n129);
and gate_103(n131,pi5,n53);
not gate_104(n132,n131);
and gate_105(n133,n130,n132);
not gate_106(n134,n133);
and gate_107(n135,n30,pi6);
not gate_108(n136,n135);
and gate_109(n137,pi0,n36);
not gate_110(n138,n137);
and gate_111(n139,n136,n138);
not gate_112(n140,n139);
and gate_113(n141,n134,n140);
and gate_114(n142,n33,n34);
not gate_115(n143,n142);
and gate_116(n144,n141,n142);
not gate_117(n145,n144);
and gate_118(n146,n35,n36);
not gate_119(n147,n146);
and gate_120(n148,n39,n146);
not gate_121(n149,n148);
and gate_122(n150,pi5,pi6);
not gate_123(n151,n150);
and gate_124(n152,n43,n150);
not gate_125(n153,n152);
and gate_126(n154,n149,n153);
not gate_127(n155,n154);
and gate_128(n156,n30,n155);
not gate_129(n157,n156);
and gate_130(n158,pi0,pi5);
and gate_131(n159,n104,n158);
not gate_132(n160,n159);
and gate_133(n161,n157,n160);
not gate_134(n162,n161);
and gate_135(n163,pi3,pi4);
not gate_136(n164,n163);
and gate_137(n165,n162,n163);
not gate_138(n166,n165);
and gate_139(n167,n145,n166);
not gate_140(n168,n167);
and gate_141(n169,n32,n168);
not gate_142(n170,n169);
and gate_143(n171,n128,n170);
not gate_144(n172,n171);
and gate_145(n173,pi1,n172);
not gate_146(n174,n173);
and gate_147(n175,pi5,n36);
not gate_148(n176,n175);
and gate_149(n177,n88,n176);
not gate_150(n178,n177);
and gate_151(n179,n36,pi7);
not gate_152(n180,n179);
and gate_153(n181,pi6,n37);
not gate_154(n182,n181);
and gate_155(n183,n180,n182);
not gate_156(n184,n183);
and gate_157(n185,pi4,n184);
not gate_158(n186,n185);
and gate_159(n187,n177,n185);
and gate_160(n188,n33,n187);
not gate_161(n189,n188);
and gate_162(n190,n98,n105);
not gate_163(n191,n190);
and gate_164(n192,pi3,n34);
not gate_165(n193,n192);
and gate_166(n194,n191,n192);
not gate_167(n195,n194);
and gate_168(n196,n189,n195);
not gate_169(n197,n196);
and gate_170(n198,n31,n197);
not gate_171(n199,n198);
and gate_172(n200,pi3,pi7);
not gate_173(n201,n200);
and gate_174(n202,n33,n37);
not gate_175(n203,n202);
and gate_176(n204,n201,n203);
not gate_177(n205,n204);
and gate_178(n206,n33,pi4);
not gate_179(n207,n206);
and gate_180(n208,n193,n207);
not gate_181(n209,n208);
and gate_182(n210,n205,n208);
and gate_183(n211,n175,n210);
not gate_184(n212,n211);
and gate_185(n213,n199,n212);
not gate_186(n214,n213);
and gate_187(n215,pi8,n214);
not gate_188(n216,n215);
and gate_189(n217,n33,pi5);
not gate_190(n218,n217);
and gate_191(n219,n33,pi7);
not gate_192(n220,n219);
and gate_193(n221,pi3,n37);
not gate_194(n222,n221);
and gate_195(n223,n220,n222);
not gate_196(n224,n223);
and gate_197(n225,pi3,pi6);
not gate_198(n226,n225);
and gate_199(n227,n33,n36);
not gate_200(n228,n227);
and gate_201(n229,n226,n228);
not gate_202(n230,n229);
and gate_203(n231,n223,n229);
and gate_204(n232,n218,n231);
and gate_205(n233,pi4,n232);
not gate_206(n234,n233);
and gate_207(n235,n176,n226);
not gate_208(n236,n235);
and gate_209(n237,pi7,n236);
not gate_210(n238,n237);
and gate_211(n239,pi3,n35);
not gate_212(n240,n239);
and gate_213(n241,n97,n239);
not gate_214(n242,n241);
and gate_215(n243,n238,n242);
not gate_216(n244,n243);
and gate_217(n245,n34,n244);
not gate_218(n246,n245);
and gate_219(n247,n234,n246);
not gate_220(n248,n247);
and gate_221(n249,n31,n38);
not gate_222(n250,n249);
and gate_223(n251,n248,n249);
not gate_224(n252,n251);
and gate_225(n253,n216,n252);
not gate_226(n254,n253);
and gate_227(n255,n32,n254);
not gate_228(n256,n255);
and gate_229(n257,pi4,pi7);
not gate_230(n258,n257);
and gate_231(n259,n40,n44);
not gate_232(n260,n259);
and gate_233(n261,n34,n260);
not gate_234(n262,n261);
and gate_235(n263,n258,n262);
not gate_236(n264,n263);
and gate_237(n265,pi5,n264);
not gate_238(n266,n265);
and gate_239(n267,n54,n82);
not gate_240(n268,n267);
and gate_241(n269,n35,n268);
not gate_242(n270,n269);
and gate_243(n271,pi4,n269);
not gate_244(n272,n271);
and gate_245(n273,n266,n272);
not gate_246(n274,n273);
and gate_247(n275,pi6,n274);
not gate_248(n276,n275);
and gate_249(n277,pi4,pi5);
not gate_250(n278,n277);
and gate_251(n279,n97,n277);
not gate_252(n280,n279);
and gate_253(n281,n276,n280);
not gate_254(n282,n281);
and gate_255(n283,pi2,n282);
not gate_256(n284,n283);
and gate_257(n285,pi4,n35);
not gate_258(n286,n285);
and gate_259(n287,n65,n285);
not gate_260(n288,n287);
and gate_261(n289,n284,n288);
not gate_262(n290,n289);
and gate_263(n291,n31,pi3);
not gate_264(n292,n291);
and gate_265(n293,n290,n291);
not gate_266(n294,n293);
and gate_267(n295,n256,n294);
not gate_268(n296,n295);
and gate_269(n297,pi0,n296);
not gate_270(n298,n297);
and gate_271(n299,n31,pi2);
not gate_272(n300,n299);
and gate_273(n301,n163,n299);
and gate_274(n302,n81,n150);
not gate_275(n303,n302);
and gate_276(n304,n301,n302);
not gate_277(n305,n304);
and gate_278(n306,n298,n305);
and gate_279(n307,n174,n306);
not gate_280(po01,n307);
and gate_281(n309,pi3,n36);
not gate_282(n310,n309);
and gate_283(n311,n52,n310);
not gate_284(n312,n311);
and gate_285(n313,n30,n31);
not gate_286(n314,n313);
and gate_287(n315,n312,n314);
not gate_288(n316,n315);
and gate_289(n317,n138,n316);
not gate_290(n318,n317);
and gate_291(n319,pi8,n318);
not gate_292(n320,n319);
and gate_293(n321,n31,n229);
not gate_294(n322,n321);
and gate_295(n323,n310,n314);
not gate_296(n324,n323);
and gate_297(n325,n322,n324);
and gate_298(n326,n38,n325);
not gate_299(n327,n326);
and gate_300(n328,n320,n327);
not gate_301(n329,n328);
and gate_302(n330,pi4,n329);
not gate_303(n331,n330);
and gate_304(n332,pi6,pi8);
not gate_305(n333,n332);
and gate_306(n334,pi3,n332);
not gate_307(n335,n334);
and gate_308(n336,n36,n38);
not gate_309(n337,n336);
and gate_310(n338,n33,n336);
not gate_311(n339,n338);
and gate_312(n340,n335,n339);
not gate_313(n341,n340);
and gate_314(n342,pi0,n341);
not gate_315(n343,n342);
and gate_316(n344,pi3,pi8);
not gate_317(n345,n344);
and gate_318(n346,n30,n38);
not gate_319(n347,n346);
and gate_320(n348,n345,n347);
not gate_321(n349,n348);
and gate_322(n350,n229,n349);
not gate_323(n351,n350);
and gate_324(n352,n343,n351);
not gate_325(n353,n352);
and gate_326(n354,pi1,n353);
not gate_327(n355,n354);
and gate_328(n356,n31,n227);
not gate_329(n357,n356);
and gate_330(n358,pi6,n38);
not gate_331(n359,n358);
and gate_332(n360,pi3,n358);
not gate_333(n361,n360);
and gate_334(n362,n357,n361);
not gate_335(n363,n362);
and gate_336(n364,pi0,n363);
not gate_337(n365,n364);
and gate_338(n366,n355,n365);
not gate_339(n367,n366);
and gate_340(n368,n34,n367);
not gate_341(n369,n368);
and gate_342(n370,n36,n310);
not gate_343(n371,n370);
and gate_344(n372,pi0,n249);
not gate_345(n373,n372);
and gate_346(n374,n371,n372);
not gate_347(n375,n374);
and gate_348(n376,n369,n375);
and gate_349(n377,n331,n376);
not gate_350(n378,n377);
and gate_351(n379,n35,n378);
not gate_352(n380,n379);
and gate_353(n381,n228,n361);
not gate_354(n382,n381);
and gate_355(n383,n31,n382);
not gate_356(n384,n383);
and gate_357(n385,n38,n230);
not gate_358(n386,n385);
and gate_359(n387,n33,pi8);
not gate_360(n388,n387);
and gate_361(n389,pi6,n387);
not gate_362(n390,n389);
and gate_363(n391,pi1,n390);
and gate_364(n392,n386,n391);
not gate_365(n393,n392);
and gate_366(n394,n384,n393);
not gate_367(n395,n394);
and gate_368(n396,pi4,n395);
not gate_369(n397,n396);
and gate_370(n398,n310,n388);
not gate_371(n399,n398);
and gate_372(n400,pi1,n399);
not gate_373(n401,n400);
and gate_374(n402,n31,n225);
not gate_375(n403,n402);
and gate_376(n404,n401,n403);
not gate_377(n405,n404);
and gate_378(n406,n34,n405);
not gate_379(n407,n406);
and gate_380(n408,n397,n407);
not gate_381(n409,n408);
and gate_382(n410,n30,n409);
not gate_383(n411,n410);
and gate_384(n412,pi4,n332);
not gate_385(n413,n412);
and gate_386(n414,pi6,n413);
not gate_387(n415,n414);
and gate_388(n416,pi1,n415);
not gate_389(n417,n416);
and gate_390(n418,n36,pi8);
not gate_391(n419,n418);
and gate_392(n420,n359,n419);
not gate_393(n421,n420);
and gate_394(n422,pi4,n36);
not gate_395(n423,n422);
and gate_396(n424,n34,pi6);
not gate_397(n425,n424);
and gate_398(n426,n423,n425);
not gate_399(n427,n426);
and gate_400(n428,n31,n426);
and gate_401(n429,n421,n428);
not gate_402(n430,n429);
and gate_403(n431,n417,n430);
not gate_404(n432,n431);
and gate_405(n433,pi3,n432);
not gate_406(n434,n433);
and gate_407(n435,n31,n34);
not gate_408(n436,n435);
and gate_409(n437,n332,n435);
not gate_410(n438,n437);
and gate_411(n439,n434,n438);
not gate_412(n440,n439);
and gate_413(n441,pi0,n440);
not gate_414(n442,n441);
and gate_415(n443,n411,n442);
not gate_416(n444,n443);
and gate_417(n445,pi5,n444);
not gate_418(n446,n445);
and gate_419(n447,n380,n446);
not gate_420(n448,n447);
and gate_421(n449,n37,n448);
not gate_422(n450,n449);
and gate_423(n451,pi4,pi8);
not gate_424(n452,n451);
and gate_425(n453,n35,n38);
not gate_426(n454,n453);
and gate_427(n455,pi5,pi8);
not gate_428(n456,n455);
and gate_429(n457,n34,n455);
not gate_430(n458,n457);
and gate_431(n459,n454,n458);
not gate_432(n460,n459);
and gate_433(n461,n452,n459);
not gate_434(n462,n461);
and gate_435(n463,n33,n462);
not gate_436(n464,n463);
and gate_437(n465,pi3,n277);
not gate_438(n466,n465);
and gate_439(n467,n464,n466);
not gate_440(n468,n467);
and gate_441(n469,pi0,n468);
not gate_442(n470,n469);
and gate_443(n471,n164,n218);
not gate_444(n472,n471);
and gate_445(n473,pi8,n472);
and gate_446(n474,n30,n473);
not gate_447(n475,n474);
and gate_448(n476,n470,n475);
not gate_449(n477,n476);
and gate_450(n478,pi6,n477);
not gate_451(n479,n478);
and gate_452(n480,pi4,n38);
not gate_453(n481,n480);
and gate_454(n482,pi3,n458);
not gate_455(n483,n482);
and gate_456(n484,n481,n483);
not gate_457(n485,n484);
and gate_458(n486,n30,n485);
not gate_459(n487,n486);
and gate_460(n488,pi3,n285);
and gate_461(n489,n347,n488);
not gate_462(n490,n489);
and gate_463(n491,n487,n490);
not gate_464(n492,n491);
and gate_465(n493,n36,n492);
not gate_466(n494,n493);
and gate_467(n495,n479,n494);
not gate_468(n496,n495);
and gate_469(n497,pi1,n496);
not gate_470(n498,n497);
and gate_471(n499,pi4,n341);
not gate_472(n500,n499);
and gate_473(n501,n36,n345);
not gate_474(n502,n501);
and gate_475(n503,n34,n502);
not gate_476(n504,n503);
and gate_477(n505,n500,n504);
not gate_478(n506,n505);
and gate_479(n507,n35,n506);
not gate_480(n508,n507);
and gate_481(n509,n34,pi5);
not gate_482(n510,n509);
and gate_483(n511,n38,n510);
not gate_484(n512,n511);
and gate_485(n513,n501,n512);
not gate_486(n514,n513);
and gate_487(n515,n508,n514);
not gate_488(n516,n515);
and gate_489(n517,pi0,n516);
not gate_490(n518,n517);
and gate_491(n519,n33,n35);
not gate_492(n520,n519);
and gate_493(n521,n33,n332);
not gate_494(n522,n521);
and gate_495(n523,n147,n522);
not gate_496(n524,n523);
and gate_497(n525,n520,n524);
and gate_498(n526,n34,n525);
not gate_499(n527,n526);
and gate_500(n528,n35,n418);
not gate_501(n529,n528);
and gate_502(n530,n36,n529);
not gate_503(n531,n530);
and gate_504(n532,n163,n531);
not gate_505(n533,n532);
and gate_506(n534,n527,n533);
not gate_507(n535,n534);
and gate_508(n536,n30,n535);
not gate_509(n537,n536);
and gate_510(n538,n518,n537);
not gate_511(n539,n538);
and gate_512(n540,n31,n539);
not gate_513(n541,n540);
and gate_514(n542,n33,n277);
not gate_515(n543,n542);
and gate_516(n544,n34,n418);
and gate_517(n545,n218,n544);
not gate_518(n546,n545);
and gate_519(n547,n543,n546);
not gate_520(n548,n547);
and gate_521(n549,pi0,n548);
not gate_522(n550,n549);
and gate_523(n551,n541,n550);
and gate_524(n552,n498,n551);
not gate_525(n553,n552);
and gate_526(n554,pi7,n553);
not gate_527(n555,n554);
and gate_528(n556,n450,n555);
not gate_529(n557,n556);
and gate_530(n558,pi2,n557);
not gate_531(n559,n558);
and gate_532(n560,pi5,n43);
not gate_533(n561,n560);
and gate_534(n562,n34,n39);
not gate_535(n563,n562);
and gate_536(n564,pi4,n62);
and gate_537(n565,n35,n564);
not gate_538(n566,n565);
and gate_539(n567,n563,n566);
and gate_540(n568,n561,n567);
not gate_541(n569,n568);
and gate_542(n570,pi6,n569);
not gate_543(n571,n570);
and gate_544(n572,n34,n453);
not gate_545(n573,n572);
and gate_546(n574,n34,n573);
not gate_547(n575,n574);
and gate_548(n576,n179,n575);
not gate_549(n577,n576);
and gate_550(n578,n571,n577);
not gate_551(n579,n578);
and gate_552(n580,n33,n579);
not gate_553(n581,n580);
and gate_554(n582,n286,n510);
not gate_555(n583,n582);
and gate_556(n584,pi6,n81);
not gate_557(n585,n584);
and gate_558(n586,n54,n585);
not gate_559(n587,n586);
and gate_560(n588,n583,n587);
not gate_561(n589,n588);
and gate_562(n590,pi5,n38);
not gate_563(n591,n590);
and gate_564(n592,n100,n591);
not gate_565(n593,n592);
and gate_566(n594,pi4,n593);
not gate_567(n595,n594);
and gate_568(n596,n34,n99);
not gate_569(n597,n596);
and gate_570(n598,n595,n597);
not gate_571(n599,n598);
and gate_572(n600,pi7,n599);
not gate_573(n601,n600);
and gate_574(n602,n81,n286);
not gate_575(n603,n602);
and gate_576(n604,n601,n603);
not gate_577(n605,n604);
and gate_578(n606,n36,n605);
not gate_579(n607,n606);
and gate_580(n608,n34,n35);
not gate_581(n609,n608);
and gate_582(n610,n43,n608);
not gate_583(n611,n610);
and gate_584(n612,n607,n611);
and gate_585(n613,n589,n612);
not gate_586(n614,n613);
and gate_587(n615,pi3,n614);
not gate_588(n616,n615);
and gate_589(n617,n36,n81);
not gate_590(n618,n617);
and gate_591(n619,n277,n617);
not gate_592(n620,n619);
and gate_593(n621,n616,n620);
and gate_594(n622,n581,n621);
not gate_595(n623,n622);
and gate_596(n624,pi0,n623);
not gate_597(n625,n624);
and gate_598(n626,pi4,pi6);
not gate_599(n627,n626);
and gate_600(n628,n81,n626);
not gate_601(n629,n628);
and gate_602(n630,n36,n53);
not gate_603(n631,n630);
and gate_604(n632,n629,n631);
not gate_605(n633,n632);
and gate_606(n634,n35,n633);
not gate_607(n635,n634);
and gate_608(n636,n34,n38);
not gate_609(n637,n636);
and gate_610(n638,n452,n637);
not gate_611(n639,n638);
and gate_612(n640,n184,n639);
not gate_613(n641,n640);
and gate_614(n642,pi4,n104);
not gate_615(n643,n642);
and gate_616(n644,n34,n97);
not gate_617(n645,n644);
and gate_618(n646,n643,n645);
not gate_619(n647,n646);
and gate_620(n648,pi8,n647);
not gate_621(n649,n648);
and gate_622(n650,n641,n649);
not gate_623(n651,n650);
and gate_624(n652,pi5,n651);
not gate_625(n653,n652);
and gate_626(n654,n635,n653);
not gate_627(n655,n654);
and gate_628(n656,pi3,n655);
not gate_629(n657,n656);
and gate_630(n658,n36,n268);
not gate_631(n659,n658);
and gate_632(n660,pi4,n658);
not gate_633(n661,n660);
and gate_634(n662,n34,pi8);
not gate_635(n663,n662);
and gate_636(n664,n481,n663);
not gate_637(n665,n664);
and gate_638(n666,pi6,n260);
not gate_639(n667,n666);
and gate_640(n668,n664,n666);
not gate_641(n669,n668);
and gate_642(n670,n661,n669);
not gate_643(n671,n670);
and gate_644(n672,n35,n671);
not gate_645(n673,n672);
and gate_646(n674,n180,n359);
and gate_647(n675,n509,n674);
not gate_648(n676,n675);
and gate_649(n677,n673,n676);
not gate_650(n678,n677);
and gate_651(n679,n33,n678);
not gate_652(n680,n679);
and gate_653(n681,n657,n680);
not gate_654(n682,n681);
and gate_655(n683,n30,n682);
not gate_656(n684,n683);
and gate_657(n685,n65,n519);
not gate_658(n686,n685);
and gate_659(n687,n684,n686);
and gate_660(n688,n625,n687);
not gate_661(n689,n688);
and gate_662(n690,pi1,n689);
not gate_663(n691,n690);
and gate_664(n692,n129,n192);
not gate_665(n693,n692);
and gate_666(n694,pi5,pi7);
not gate_667(n695,n694);
and gate_668(n696,n33,n694);
and gate_669(n697,n665,n696);
not gate_670(n698,n697);
and gate_671(n699,n693,n698);
and gate_672(n700,n53,n146);
not gate_673(n701,n700);
and gate_674(n702,n303,n701);
not gate_675(n703,n702);
and gate_676(n704,n34,n703);
not gate_677(n705,n704);
and gate_678(n706,pi5,n37);
not gate_679(n707,n706);
and gate_680(n708,n35,n39);
not gate_681(n709,n708);
and gate_682(n710,n707,n709);
not gate_683(n711,n710);
and gate_684(n712,pi6,n711);
not gate_685(n713,n712);
and gate_686(n714,n418,n695);
not gate_687(n715,n714);
and gate_688(n716,n713,n715);
not gate_689(n717,n716);
and gate_690(n718,pi4,n717);
not gate_691(n719,n718);
and gate_692(n720,n705,n719);
not gate_693(n721,n720);
and gate_694(n722,pi3,n721);
not gate_695(n723,n722);
and gate_696(n724,n43,n175);
not gate_697(n725,n724);
and gate_698(n726,pi5,n48);
not gate_699(n727,n726);
and gate_700(n728,n35,n332);
not gate_701(n729,n728);
and gate_702(n730,n727,n729);
not gate_703(n731,n730);
and gate_704(n732,n206,n731);
not gate_705(n733,n732);
and gate_706(n734,n725,n733);
and gate_707(n735,n723,n734);
and gate_708(n736,n699,n735);
not gate_709(n737,n736);
and gate_710(n738,n31,n737);
not gate_711(n739,n738);
and gate_712(n740,n107,n707);
not gate_713(n741,n740);
and gate_714(n742,n34,n741);
not gate_715(n743,n742);
and gate_716(n744,pi4,n146);
not gate_717(n745,n744);
and gate_718(n746,n743,n745);
not gate_719(n747,n746);
and gate_720(n748,n33,n38);
not gate_721(n749,n748);
and gate_722(n750,n747,n748);
not gate_723(n751,n750);
and gate_724(n752,n739,n751);
not gate_725(n753,n752);
and gate_726(n754,pi0,n753);
not gate_727(n755,n754);
and gate_728(n756,n691,n755);
not gate_729(n757,n756);
and gate_730(n758,n32,n757);
not gate_731(n759,n758);
and gate_732(n760,n34,n179);
not gate_733(n761,n760);
and gate_734(n762,pi4,n706);
not gate_735(n763,n762);
and gate_736(n764,n761,n763);
not gate_737(n765,n764);
and gate_738(n766,pi0,n765);
not gate_739(n767,n766);
and gate_740(n768,n30,pi4);
not gate_741(n769,n768);
and gate_742(n770,n35,n181);
and gate_743(n771,n768,n770);
not gate_744(n772,n771);
and gate_745(n773,n767,n772);
not gate_746(n774,n773);
and gate_747(n775,pi3,n774);
not gate_748(n776,n775);
and gate_749(n777,n30,n142);
and gate_750(n778,n106,n777);
not gate_751(n779,n778);
and gate_752(n780,n776,n779);
not gate_753(n781,n780);
and gate_754(n782,n38,n781);
not gate_755(n783,n782);
and gate_756(n784,n34,n36);
not gate_757(n785,n784);
and gate_758(n786,n33,n784);
not gate_759(n787,n786);
and gate_760(n788,n226,n787);
not gate_761(n789,n788);
and gate_762(n790,pi5,n39);
not gate_763(n791,n790);
and gate_764(n792,n789,n790);
and gate_765(n793,pi0,n792);
not gate_766(n794,n793);
and gate_767(n795,n783,n794);
not gate_768(n796,n795);
and gate_769(n797,pi1,n796);
not gate_770(n798,n797);
and gate_771(n799,n31,n33);
not gate_772(n800,n799);
and gate_773(n801,pi0,n799);
and gate_774(n802,n34,n181);
not gate_775(n803,n802);
and gate_776(n804,n456,n802);
and gate_777(n805,n801,n804);
not gate_778(n806,n805);
and gate_779(n807,n798,n806);
and gate_780(n808,n759,n807);
and gate_781(n809,n559,n808);
not gate_782(po02,n809);
and gate_783(n811,pi4,n99);
not gate_784(n812,n811);
and gate_785(n813,n34,n590);
not gate_786(n814,n813);
and gate_787(n815,n812,n814);
not gate_788(n816,n815);
and gate_789(n817,n32,pi3);
not gate_790(n818,n817);
and gate_791(n819,pi2,n33);
not gate_792(n820,n819);
and gate_793(n821,n818,n820);
not gate_794(n822,n821);
and gate_795(n823,n97,n822);
and gate_796(n824,pi1,n823);
not gate_797(n825,n824);
and gate_798(n826,n33,n104);
and gate_799(n827,n299,n826);
not gate_800(n828,n827);
and gate_801(n829,n825,n828);
not gate_802(n830,n829);
and gate_803(n831,n816,n830);
not gate_804(n832,n831);
and gate_805(n833,n585,n631);
not gate_806(n834,n833);
and gate_807(n835,n31,n834);
not gate_808(n836,n835);
and gate_809(n837,pi6,n268);
not gate_810(n838,n837);
and gate_811(n839,n98,n838);
not gate_812(n840,n839);
and gate_813(n841,pi1,n840);
not gate_814(n842,n841);
and gate_815(n843,n836,n842);
not gate_816(n844,n843);
and gate_817(n845,n35,n844);
not gate_818(n846,n845);
and gate_819(n847,n82,n631);
and gate_820(n848,n667,n847);
not gate_821(n849,n848);
and gate_822(n850,pi1,n849);
not gate_823(n851,n850);
and gate_824(n852,n31,n37);
not gate_825(n853,n852);
and gate_826(n854,n358,n852);
not gate_827(n855,n854);
and gate_828(n856,n851,n855);
not gate_829(n857,n856);
and gate_830(n858,pi5,n857);
not gate_831(n859,n858);
and gate_832(n860,n846,n859);
not gate_833(n861,n860);
and gate_834(n862,pi4,n861);
not gate_835(n863,n862);
and gate_836(n864,n36,n100);
and gate_837(n865,n54,n864);
not gate_838(n866,n865);
and gate_839(n867,n107,n866);
not gate_840(n868,n867);
and gate_841(n869,pi1,n34);
and gate_842(n870,n868,n869);
not gate_843(n871,n870);
and gate_844(n872,n863,n871);
not gate_845(n873,n872);
and gate_846(n874,pi3,n873);
not gate_847(n875,n874);
and gate_848(n876,n43,n423);
not gate_849(n877,n876);
and gate_850(n878,n42,n877);
not gate_851(n879,n878);
and gate_852(n880,n35,n879);
not gate_853(n881,n880);
and gate_854(n882,n36,n40);
not gate_855(n883,n882);
and gate_856(n884,n34,pi7);
not gate_857(n885,n884);
and gate_858(n886,pi4,n37);
not gate_859(n887,n886);
and gate_860(n888,n885,n887);
not gate_861(n889,n888);
and gate_862(n890,n82,n889);
not gate_863(n891,n890);
and gate_864(n892,n883,n891);
and gate_865(n893,pi5,n892);
not gate_866(n894,n893);
and gate_867(n895,n881,n894);
not gate_868(n896,n895);
and gate_869(n897,pi1,n33);
not gate_870(n898,n897);
and gate_871(n899,n896,n897);
not gate_872(n900,n899);
and gate_873(n901,n875,n900);
not gate_874(n902,n901);
and gate_875(n903,pi2,n902);
not gate_876(n904,n903);
and gate_877(n905,pi6,n39);
not gate_878(n906,n905);
and gate_879(n907,n32,n34);
not gate_880(n908,n907);
and gate_881(n909,n905,n907);
not gate_882(n910,n909);
and gate_883(n911,n43,n422);
not gate_884(n912,n911);
and gate_885(n913,n910,n912);
not gate_886(n914,n913);
and gate_887(n915,n33,n914);
not gate_888(n916,n915);
and gate_889(n917,n180,n803);
not gate_890(n918,n917);
and gate_891(n919,pi8,n918);
and gate_892(n920,n817,n919);
not gate_893(n921,n920);
and gate_894(n922,n916,n921);
not gate_895(n923,n922);
and gate_896(n924,pi5,n923);
not gate_897(n925,n924);
and gate_898(n926,n99,n142);
not gate_899(n927,n926);
and gate_900(n928,pi3,n480);
not gate_901(n929,n928);
and gate_902(n930,n927,n929);
and gate_903(n931,n35,n358);
and gate_904(n932,n33,n931);
not gate_905(n933,n932);
and gate_906(n934,n930,n933);
not gate_907(n935,n934);
and gate_908(n936,pi7,n935);
not gate_909(n937,n936);
and gate_910(n938,n192,n528);
not gate_911(n939,n938);
and gate_912(n940,n937,n939);
not gate_913(n941,n940);
and gate_914(n942,n32,n941);
not gate_915(n943,n942);
and gate_916(n944,n925,n943);
not gate_917(n945,n944);
and gate_918(n946,pi1,n945);
not gate_919(n947,n946);
and gate_920(n948,n904,n947);
and gate_921(n949,n832,n948);
not gate_922(n950,n949);
and gate_923(n951,n30,n950);
not gate_924(n952,n951);
and gate_925(n953,pi1,pi3);
not gate_926(n954,n953);
and gate_927(n955,n790,n953);
not gate_928(n956,n955);
and gate_929(n957,n35,n43);
not gate_930(n958,n957);
and gate_931(n959,n799,n957);
not gate_932(n960,n959);
and gate_933(n961,n956,n960);
not gate_934(n962,n961);
and gate_935(n963,n36,n962);
not gate_936(n964,n963);
and gate_937(n965,n31,pi8);
not gate_938(n966,n965);
and gate_939(n967,n454,n966);
not gate_940(n968,n967);
and gate_941(n969,pi1,pi7);
not gate_942(n970,n969);
and gate_943(n971,n707,n970);
not gate_944(n972,n971);
and gate_945(n973,n968,n972);
and gate_946(n974,n33,n973);
not gate_947(n975,n974);
and gate_948(n976,n853,n970);
not gate_949(n977,n976);
and gate_950(n978,n35,n977);
not gate_951(n979,n978);
and gate_952(n980,n31,pi5);
not gate_953(n981,n980);
and gate_954(n982,n53,n980);
not gate_955(n983,n982);
and gate_956(n984,n979,n983);
not gate_957(n985,n984);
and gate_958(n986,pi3,n985);
not gate_959(n987,n986);
and gate_960(n988,n975,n987);
not gate_961(n989,n988);
and gate_962(n990,pi6,n989);
not gate_963(n991,n990);
and gate_964(n992,n964,n991);
not gate_965(n993,n992);
and gate_966(n994,pi2,n993);
not gate_967(n995,n994);
and gate_968(n996,pi5,n104);
not gate_969(n997,n996);
and gate_970(n998,n35,n97);
not gate_971(n999,n998);
and gate_972(n1000,n997,n999);
not gate_973(n1001,n1000);
and gate_974(n1002,n33,n1001);
not gate_975(n1003,n1002);
and gate_976(n1004,n35,pi7);
not gate_977(n1005,n1004);
and gate_978(n1006,n707,n1005);
not gate_979(n1007,n1006);
and gate_980(n1008,pi6,n1007);
not gate_981(n1009,n1008);
and gate_982(n1010,n1003,n1009);
not gate_983(n1011,n1010);
and gate_984(n1012,pi8,n1011);
not gate_985(n1013,n1012);
and gate_986(n1014,pi8,n147);
not gate_987(n1015,n1014);
and gate_988(n1016,n1006,n1015);
and gate_989(n1017,pi3,n1016);
not gate_990(n1018,n1017);
and gate_991(n1019,n1013,n1018);
not gate_992(n1020,n1019);
and gate_993(n1021,pi1,n1020);
not gate_994(n1022,n1021);
and gate_995(n1023,n44,n906);
not gate_996(n1024,n1023);
and gate_997(n1025,pi3,n39);
not gate_998(n1026,n1025);
and gate_999(n1027,n311,n1026);
not gate_1000(n1028,n1027);
and gate_1001(n1029,n1024,n1028);
and gate_1002(n1030,pi5,n1029);
not gate_1003(n1031,n1030);
and gate_1004(n1032,n335,n749);
not gate_1005(n1033,n1032);
and gate_1006(n1034,pi7,n1033);
not gate_1007(n1035,n1034);
and gate_1008(n1036,n618,n1035);
not gate_1009(n1037,n1036);
and gate_1010(n1038,n35,n1037);
not gate_1011(n1039,n1038);
and gate_1012(n1040,n1031,n1039);
not gate_1013(n1041,n1040);
and gate_1014(n1042,n31,n1041);
not gate_1015(n1043,n1042);
and gate_1016(n1044,n1022,n1043);
not gate_1017(n1045,n1044);
and gate_1018(n1046,n32,n1045);
not gate_1019(n1047,n1046);
and gate_1020(n1048,pi1,n36);
not gate_1021(n1049,n1048);
and gate_1022(n1050,n31,n176);
not gate_1023(n1051,n1050);
and gate_1024(n1052,n1049,n1051);
and gate_1025(n1053,n81,n1052);
and gate_1026(n1054,n33,n1053);
not gate_1027(n1055,n1054);
and gate_1028(n1056,n1047,n1055);
and gate_1029(n1057,n995,n1056);
not gate_1030(n1058,n1057);
and gate_1031(n1059,pi4,n1058);
not gate_1032(n1060,n1059);
and gate_1033(n1061,n706,n817);
not gate_1034(n1062,n1061);
and gate_1035(n1063,pi2,n35);
not gate_1036(n1064,n1063);
and gate_1037(n1065,pi3,n1063);
not gate_1038(n1066,n1065);
and gate_1039(n1067,pi7,n1066);
and gate_1040(n1068,n115,n520);
not gate_1041(n1069,n1068);
and gate_1042(n1070,n32,n1069);
not gate_1043(n1071,n1070);
and gate_1044(n1072,n1067,n1071);
not gate_1045(n1073,n1072);
and gate_1046(n1074,n1062,n1073);
not gate_1047(n1075,n1074);
and gate_1048(n1076,n31,n1075);
not gate_1049(n1077,n1076);
and gate_1050(n1078,n35,n37);
not gate_1051(n1079,n1078);
and gate_1052(n1080,n33,n1079);
not gate_1053(n1081,n1080);
and gate_1054(n1082,pi2,n1081);
not gate_1055(n1083,n1082);
and gate_1056(n1084,n32,pi5);
not gate_1057(n1085,n1084);
and gate_1058(n1086,n224,n1084);
not gate_1059(n1087,n1086);
and gate_1060(n1088,n1083,n1087);
not gate_1061(n1089,n1088);
and gate_1062(n1090,pi1,n1089);
not gate_1063(n1091,n1090);
and gate_1064(n1092,n1077,n1091);
not gate_1065(n1093,n1092);
and gate_1066(n1094,pi6,n1093);
not gate_1067(n1095,n1094);
and gate_1068(n1096,n1064,n1085);
not gate_1069(n1097,n1096);
and gate_1070(n1098,pi1,n1097);
not gate_1071(n1099,n1098);
and gate_1072(n1100,n32,n35);
not gate_1073(n1101,n1100);
and gate_1074(n1102,n31,n1100);
not gate_1075(n1103,n1102);
and gate_1076(n1104,n1099,n1103);
not gate_1077(n1105,n1104);
and gate_1078(n1106,pi3,n1105);
not gate_1079(n1107,n1106);
and gate_1080(n1108,pi1,pi5);
not gate_1081(n1109,n1108);
and gate_1082(n1110,n818,n1064);
and gate_1083(n1111,n1109,n1110);
not gate_1084(n1112,n1111);
and gate_1085(n1113,n1107,n1112);
not gate_1086(n1114,n1113);
and gate_1087(n1115,n37,n1114);
not gate_1088(n1116,n1115);
and gate_1089(n1117,n299,n1004);
not gate_1090(n1118,n1117);
and gate_1091(n1119,n1116,n1118);
not gate_1092(n1120,n1119);
and gate_1093(n1121,n36,n1120);
not gate_1094(n1122,n1121);
and gate_1095(n1123,n1095,n1122);
not gate_1096(n1124,n1123);
and gate_1097(n1125,n38,n1124);
not gate_1098(n1126,n1125);
and gate_1099(n1127,n695,n1079);
not gate_1100(n1128,n1127);
and gate_1101(n1129,n31,n1128);
not gate_1102(n1130,n1129);
and gate_1103(n1131,pi1,n1004);
not gate_1104(n1132,n1131);
and gate_1105(n1133,n1130,n1132);
not gate_1106(n1134,n1133);
and gate_1107(n1135,pi3,n1134);
not gate_1108(n1136,n1135);
and gate_1109(n1137,pi1,pi2);
not gate_1110(n1138,n1137);
and gate_1111(n1139,n217,n1137);
not gate_1112(n1140,n1139);
and gate_1113(n1141,n1136,n1140);
not gate_1114(n1142,n1141);
and gate_1115(n1143,pi8,n1142);
not gate_1116(n1144,n1143);
and gate_1117(n1145,pi1,n32);
not gate_1118(n1146,n1145);
and gate_1119(n1147,n33,n1004);
and gate_1120(n1148,n1145,n1147);
not gate_1121(n1149,n1148);
and gate_1122(n1150,n1144,n1149);
not gate_1123(n1151,n1150);
and gate_1124(n1152,pi6,n1151);
not gate_1125(n1153,n1152);
and gate_1126(n1154,n32,n33);
and gate_1127(n1155,n31,n36);
not gate_1128(n1156,n1155);
and gate_1129(n1157,n39,n1155);
not gate_1130(n1158,n1157);
and gate_1131(n1159,n1154,n1157);
not gate_1132(n1160,n1159);
and gate_1133(n1161,n1153,n1160);
and gate_1134(n1162,n1126,n1161);
not gate_1135(n1163,n1162);
and gate_1136(n1164,n34,n1163);
not gate_1137(n1165,n1164);
and gate_1138(n1166,n31,n819);
and gate_1139(n1167,pi5,n97);
not gate_1140(n1168,n1167);
and gate_1141(n1169,n1166,n1167);
not gate_1142(n1170,n1169);
and gate_1143(n1171,n1165,n1170);
and gate_1144(n1172,n1060,n1171);
not gate_1145(n1173,n1172);
and gate_1146(n1174,pi0,n1173);
not gate_1147(n1175,n1174);
and gate_1148(n1176,n32,pi7);
not gate_1149(n1177,n1176);
and gate_1150(n1178,pi2,n37);
not gate_1151(n1179,n1178);
and gate_1152(n1180,n1177,n1179);
not gate_1153(n1181,n1180);
and gate_1154(n1182,n32,pi4);
not gate_1155(n1183,n1182);
and gate_1156(n1184,pi2,n34);
not gate_1157(n1185,n1184);
and gate_1158(n1186,n1183,n1185);
not gate_1159(n1187,n1186);
and gate_1160(n1188,n38,n1187);
and gate_1161(n1189,n1180,n1188);
and gate_1162(n1190,n897,n1189);
not gate_1163(n1191,n1190);
and gate_1164(n1192,pi2,pi3);
not gate_1165(n1193,n1192);
and gate_1166(n1194,n31,n39);
not gate_1167(n1195,n1194);
and gate_1168(n1196,n1192,n1194);
not gate_1169(n1197,n1196);
and gate_1170(n1198,n1191,n1197);
not gate_1171(n1199,n1198);
and gate_1172(n1200,pi5,n1199);
not gate_1173(n1201,n1200);
and gate_1174(n1202,n292,n898);
not gate_1175(n1203,n1202);
and gate_1176(n1204,n224,n1203);
and gate_1177(n1205,n596,n1204);
and gate_1178(n1206,pi2,n1205);
not gate_1179(n1207,n1206);
and gate_1180(n1208,n1201,n1207);
not gate_1181(n1209,n1208);
and gate_1182(n1210,n36,n1209);
not gate_1183(n1211,n1210);
and gate_1184(n1212,n1175,n1211);
and gate_1185(n1213,n952,n1212);
not gate_1186(po03,n1213);
and gate_1187(n1215,n30,n32);
and gate_1188(n1216,pi5,n418);
not gate_1189(n1217,n1216);
and gate_1190(n1218,n1215,n1216);
not gate_1191(n1219,n1218);
and gate_1192(n1220,pi2,n99);
not gate_1193(n1221,n1220);
and gate_1194(n1222,n32,n590);
not gate_1195(n1223,n1222);
and gate_1196(n1224,pi0,n1222);
not gate_1197(n1225,n1224);
and gate_1198(n1226,n1221,n1225);
not gate_1199(n1227,n1226);
and gate_1200(n1228,pi6,n1227);
not gate_1201(n1229,n1228);
and gate_1202(n1230,n1219,n1229);
not gate_1203(n1231,n1230);
and gate_1204(n1232,pi3,n1231);
not gate_1205(n1233,n1232);
and gate_1206(n1234,pi0,n819);
and gate_1207(n1235,n931,n1234);
not gate_1208(n1236,n1235);
and gate_1209(n1237,n1233,n1236);
not gate_1210(n1238,n1237);
and gate_1211(n1239,pi1,n1238);
not gate_1212(n1240,n1239);
and gate_1213(n1241,n31,n32);
not gate_1214(n1242,n1241);
and gate_1215(n1243,pi0,n1241);
and gate_1216(n1244,n217,n336);
and gate_1217(n1245,n1243,n1244);
not gate_1218(n1246,n1245);
and gate_1219(n1247,n1240,n1246);
not gate_1220(n1248,n1247);
and gate_1221(n1249,pi4,n1248);
not gate_1222(n1250,n1249);
and gate_1223(n1251,n300,n1146);
not gate_1224(n1252,n1251);
and gate_1225(n1253,n218,n240);
not gate_1226(n1254,n1253);
and gate_1227(n1255,n1096,n1253);
and gate_1228(n1256,n1252,n1255);
and gate_1229(n1257,pi0,n1256);
not gate_1230(n1258,n1257);
and gate_1231(n1259,n30,n299);
and gate_1232(n1260,n217,n1259);
not gate_1233(n1261,n1260);
and gate_1234(n1262,n1258,n1261);
not gate_1235(n1263,n1262);
and gate_1236(n1264,n34,n332);
not gate_1237(n1265,n1264);
and gate_1238(n1266,n1263,n1264);
not gate_1239(n1267,n1266);
and gate_1240(n1268,n1250,n1267);
and gate_1241(n1269,n34,n81);
not gate_1242(n1270,n1269);
and gate_1243(n1271,n1145,n1269);
not gate_1244(n1272,n1271);
and gate_1245(n1273,pi4,n53);
not gate_1246(n1274,n1273);
and gate_1247(n1275,n299,n1273);
not gate_1248(n1276,n1275);
and gate_1249(n1277,n1272,n1276);
not gate_1250(n1278,n1277);
and gate_1251(n1279,n1069,n1278);
not gate_1252(n1280,n1279);
and gate_1253(n1281,n481,n563);
not gate_1254(n1282,n1281);
and gate_1255(n1283,pi3,n1282);
not gate_1256(n1284,n1283);
and gate_1257(n1285,pi4,n81);
not gate_1258(n1286,n1285);
and gate_1259(n1287,n34,n53);
not gate_1260(n1288,n1287);
and gate_1261(n1289,n1286,n1288);
not gate_1262(n1290,n1289);
and gate_1263(n1291,n33,n1290);
not gate_1264(n1292,n1291);
and gate_1265(n1293,n1284,n1292);
not gate_1266(n1294,n1293);
and gate_1267(n1295,n32,n1294);
not gate_1268(n1296,n1295);
and gate_1269(n1297,n53,n163);
not gate_1270(n1298,n1297);
and gate_1271(n1299,pi3,n38);
not gate_1272(n1300,n1299);
and gate_1273(n1301,n37,n1299);
not gate_1274(n1302,n1301);
and gate_1275(n1303,n34,n1302);
and gate_1276(n1304,n33,n268);
not gate_1277(n1305,n1304);
and gate_1278(n1306,n1303,n1305);
not gate_1279(n1307,n1306);
and gate_1280(n1308,n1298,n1307);
not gate_1281(n1309,n1308);
and gate_1282(n1310,pi2,n1309);
not gate_1283(n1311,n1310);
and gate_1284(n1312,n1296,n1311);
not gate_1285(n1313,n1312);
and gate_1286(n1314,n35,n1313);
not gate_1287(n1315,n1314);
and gate_1288(n1316,pi2,n163);
not gate_1289(n1317,n1316);
and gate_1290(n1318,n32,n142);
not gate_1291(n1319,n1318);
and gate_1292(n1320,n1317,n1319);
not gate_1293(n1321,n1320);
and gate_1294(n1322,n260,n1321);
not gate_1295(n1323,n1322);
and gate_1296(n1324,n34,n37);
not gate_1297(n1325,n1324);
and gate_1298(n1326,pi4,n268);
not gate_1299(n1327,n1326);
and gate_1300(n1328,n1325,n1327);
not gate_1301(n1329,n1328);
and gate_1302(n1330,n819,n1329);
not gate_1303(n1331,n1330);
and gate_1304(n1332,n1323,n1331);
not gate_1305(n1333,n1332);
and gate_1306(n1334,pi5,n1333);
not gate_1307(n1335,n1334);
and gate_1308(n1336,n562,n1192);
not gate_1309(n1337,n1336);
and gate_1310(n1338,n1335,n1337);
and gate_1311(n1339,n1315,n1338);
not gate_1312(n1340,n1339);
and gate_1313(n1341,pi1,n1340);
not gate_1314(n1342,n1341);
and gate_1315(n1343,n1280,n1342);
not gate_1316(n1344,n1343);
and gate_1317(n1345,n30,n1344);
not gate_1318(n1346,n1345);
and gate_1319(n1347,pi1,n1182);
not gate_1320(n1348,n1347);
and gate_1321(n1349,n799,n1186);
not gate_1322(n1350,n1349);
and gate_1323(n1351,n1348,n1350);
not gate_1324(n1352,n1351);
and gate_1325(n1353,pi8,n1352);
not gate_1326(n1354,n1353);
and gate_1327(n1355,n345,n749);
not gate_1328(n1356,n1355);
and gate_1329(n1357,pi2,n1356);
not gate_1330(n1358,n1357);
and gate_1331(n1359,n32,n1299);
not gate_1332(n1360,n1359);
and gate_1333(n1361,n1358,n1360);
not gate_1334(n1362,n1361);
and gate_1335(n1363,pi1,pi4);
not gate_1336(n1364,n1363);
and gate_1337(n1365,n436,n1364);
not gate_1338(n1366,n1365);
and gate_1339(n1367,n1362,n1365);
not gate_1340(n1368,n1367);
and gate_1341(n1369,n1354,n1368);
not gate_1342(n1370,n1369);
and gate_1343(n1371,n37,n1370);
not gate_1344(n1372,n1371);
and gate_1345(n1373,n800,n1356);
not gate_1346(n1374,n1373);
and gate_1347(n1375,n37,n954);
not gate_1348(n1376,n1375);
and gate_1349(n1377,n1374,n1376);
and gate_1350(n1378,pi2,n1377);
not gate_1351(n1379,n1378);
and gate_1352(n1380,pi3,n53);
and gate_1353(n1381,n1241,n1380);
not gate_1354(n1382,n1381);
and gate_1355(n1383,n1379,n1382);
not gate_1356(n1384,n1383);
and gate_1357(n1385,n34,n1384);
not gate_1358(n1386,n1385);
and gate_1359(n1387,n33,n257);
and gate_1360(n1388,n32,n1387);
not gate_1361(n1389,n1388);
and gate_1362(n1390,n1386,n1389);
and gate_1363(n1391,n1372,n1390);
not gate_1364(n1392,n1391);
and gate_1365(n1393,pi5,n1392);
not gate_1366(n1394,n1393);
and gate_1367(n1395,pi2,n889);
not gate_1368(n1396,n1395);
and gate_1369(n1397,n32,n257);
not gate_1370(n1398,n1397);
and gate_1371(n1399,n1396,n1398);
not gate_1372(n1400,n1399);
and gate_1373(n1401,n38,n1400);
not gate_1374(n1402,n1401);
and gate_1375(n1403,n81,n907);
not gate_1376(n1404,n1403);
and gate_1377(n1405,n1402,n1404);
not gate_1378(n1406,n1405);
and gate_1379(n1407,pi3,n1406);
not gate_1380(n1408,n1407);
and gate_1381(n1409,n38,n1179);
not gate_1382(n1410,n1409);
and gate_1383(n1411,n888,n1410);
and gate_1384(n1412,n33,n1411);
not gate_1385(n1413,n1412);
and gate_1386(n1414,n1408,n1413);
not gate_1387(n1415,n1414);
and gate_1388(n1416,n31,n1415);
not gate_1389(n1417,n1416);
and gate_1390(n1418,pi2,n665);
not gate_1391(n1419,n1418);
and gate_1392(n1420,n908,n1419);
not gate_1393(n1421,n1420);
and gate_1394(n1422,pi7,n1421);
not gate_1395(n1423,n1422);
and gate_1396(n1424,n81,n1182);
not gate_1397(n1425,n1424);
and gate_1398(n1426,n1423,n1425);
not gate_1399(n1427,n1426);
and gate_1400(n1428,pi3,n1427);
not gate_1401(n1429,n1428);
and gate_1402(n1430,pi4,n43);
not gate_1403(n1431,n1430);
and gate_1404(n1432,n1154,n1430);
not gate_1405(n1433,n1432);
and gate_1406(n1434,n1429,n1433);
not gate_1407(n1435,n1434);
and gate_1408(n1436,pi1,n1435);
not gate_1409(n1437,n1436);
and gate_1410(n1438,n1417,n1437);
not gate_1411(n1439,n1438);
and gate_1412(n1440,n35,n1439);
not gate_1413(n1441,n1440);
and gate_1414(n1442,n1394,n1441);
not gate_1415(n1443,n1442);
and gate_1416(n1444,pi0,n1443);
not gate_1417(n1445,n1444);
and gate_1418(n1446,n1346,n1445);
not gate_1419(n1447,n1446);
and gate_1420(n1448,pi6,n1447);
not gate_1421(n1449,n1448);
and gate_1422(n1450,n1078,n1145);
not gate_1423(n1451,n1450);
and gate_1424(n1452,pi2,n694);
not gate_1425(n1453,n1452);
and gate_1426(n1454,n31,n1452);
not gate_1427(n1455,n1454);
and gate_1428(n1456,n1451,n1455);
and gate_1429(n1457,n590,n1181);
and gate_1430(n1458,pi1,n1457);
not gate_1431(n1459,n1458);
and gate_1432(n1460,n129,n299);
not gate_1433(n1461,n1460);
and gate_1434(n1462,n1459,n1461);
and gate_1435(n1463,n1456,n1462);
not gate_1436(n1464,n1463);
and gate_1437(n1465,pi4,n1464);
not gate_1438(n1466,n1465);
and gate_1439(n1467,n39,n1145);
not gate_1440(n1468,n1467);
and gate_1441(n1469,n43,n1242);
not gate_1442(n1470,n1469);
and gate_1443(n1471,n1468,n1470);
not gate_1444(n1472,n1471);
and gate_1445(n1473,n35,n1472);
not gate_1446(n1474,n1473);
and gate_1447(n1475,pi2,n53);
not gate_1448(n1476,n1475);
and gate_1449(n1477,n1474,n1476);
not gate_1450(n1478,n1477);
and gate_1451(n1479,n34,n1478);
not gate_1452(n1480,n1479);
and gate_1453(n1481,n1466,n1480);
not gate_1454(n1482,n1481);
and gate_1455(n1483,n30,n1482);
not gate_1456(n1484,n1483);
and gate_1457(n1485,n662,n1109);
and gate_1458(n1486,pi2,n1485);
not gate_1459(n1487,n1486);
and gate_1460(n1488,n32,n38);
not gate_1461(n1489,n1488);
and gate_1462(n1490,n278,n609);
not gate_1463(n1491,n1490);
and gate_1464(n1492,n31,n1491);
not gate_1465(n1493,n1492);
and gate_1466(n1494,pi1,n285);
not gate_1467(n1495,n1494);
and gate_1468(n1496,n1109,n1495);
and gate_1469(n1497,n1493,n1496);
not gate_1470(n1498,n1497);
and gate_1471(n1499,n1488,n1498);
not gate_1472(n1500,n1499);
and gate_1473(n1501,n1487,n1500);
not gate_1474(n1502,n1501);
and gate_1475(n1503,n37,n1502);
not gate_1476(n1504,n1503);
and gate_1477(n1505,n32,pi8);
not gate_1478(n1506,n1505);
and gate_1479(n1507,pi2,n480);
not gate_1480(n1508,n1507);
and gate_1481(n1509,n1506,n1508);
not gate_1482(n1510,n1509);
and gate_1483(n1511,n31,n1510);
not gate_1484(n1512,n1511);
and gate_1485(n1513,n451,n1137);
not gate_1486(n1514,n1513);
and gate_1487(n1515,n1512,n1514);
not gate_1488(n1516,n1515);
and gate_1489(n1517,n694,n1516);
not gate_1490(n1518,n1517);
and gate_1491(n1519,n1504,n1518);
not gate_1492(n1520,n1519);
and gate_1493(n1521,pi0,n1520);
not gate_1494(n1522,n1521);
and gate_1495(n1523,n1484,n1522);
not gate_1496(n1524,n1523);
and gate_1497(n1525,pi3,n1524);
not gate_1498(n1526,n1525);
and gate_1499(n1527,pi1,n38);
not gate_1500(n1528,n1527);
and gate_1501(n1529,n35,n481);
not gate_1502(n1530,n1529);
and gate_1503(n1531,n1528,n1530);
and gate_1504(n1532,pi0,n1531);
not gate_1505(n1533,n1532);
and gate_1506(n1534,pi1,pi8);
not gate_1507(n1535,n1534);
and gate_1508(n1536,n30,n1534);
not gate_1509(n1537,n1536);
and gate_1510(n1538,pi8,n1537);
not gate_1511(n1539,n1538);
and gate_1512(n1540,n277,n1539);
not gate_1513(n1541,n1540);
and gate_1514(n1542,pi1,n35);
not gate_1515(n1543,n1542);
and gate_1516(n1544,n30,n1542);
and gate_1517(n1545,n452,n1544);
not gate_1518(n1546,n1545);
and gate_1519(n1547,n1541,n1546);
and gate_1520(n1548,n1533,n1547);
not gate_1521(n1549,n1548);
and gate_1522(n1550,pi2,n1549);
not gate_1523(n1551,n1550);
and gate_1524(n1552,n30,n34);
not gate_1525(n1553,n1552);
and gate_1526(n1554,n638,n1553);
and gate_1527(n1555,n250,n1554);
and gate_1528(n1556,pi5,n1555);
not gate_1529(n1557,n1556);
and gate_1530(n1558,n608,n1535);
and gate_1531(n1559,pi0,n1558);
not gate_1532(n1560,n1559);
and gate_1533(n1561,n1557,n1560);
not gate_1534(n1562,n1561);
and gate_1535(n1563,n32,n1562);
not gate_1536(n1564,n1563);
and gate_1537(n1565,n1551,n1564);
not gate_1538(n1566,n1565);
and gate_1539(n1567,n37,n1566);
not gate_1540(n1568,n1567);
and gate_1541(n1569,n32,n454);
not gate_1542(n1570,n1569);
and gate_1543(n1571,n30,n1570);
not gate_1544(n1572,n1571);
and gate_1545(n1573,n1225,n1572);
not gate_1546(n1574,n1573);
and gate_1547(n1575,pi1,n1574);
not gate_1548(n1576,n1575);
and gate_1549(n1577,pi2,pi5);
not gate_1550(n1578,n1577);
and gate_1551(n1579,n965,n1578);
and gate_1552(n1580,pi0,n1579);
not gate_1553(n1581,n1580);
and gate_1554(n1582,n1576,n1581);
not gate_1555(n1583,n1582);
and gate_1556(n1584,n34,n1583);
not gate_1557(n1585,n1584);
and gate_1558(n1586,n30,pi1);
not gate_1559(n1587,n1586);
and gate_1560(n1588,n1220,n1586);
not gate_1561(n1589,n1588);
and gate_1562(n1590,n1585,n1589);
not gate_1563(n1591,n1590);
and gate_1564(n1592,pi7,n1591);
not gate_1565(n1593,n1592);
and gate_1566(n1594,n572,n1243);
not gate_1567(n1595,n1594);
and gate_1568(n1596,n1593,n1595);
and gate_1569(n1597,n1568,n1596);
not gate_1570(n1598,n1597);
and gate_1571(n1599,n33,n1598);
not gate_1572(n1600,n1599);
and gate_1573(n1601,n590,n1363);
not gate_1574(n1602,n1601);
and gate_1575(n1603,n597,n1602);
not gate_1576(n1604,n1603);
and gate_1577(n1605,pi2,n1604);
not gate_1578(n1606,n1605);
and gate_1579(n1607,n592,n665);
and gate_1580(n1608,n1145,n1607);
not gate_1581(n1609,n1608);
and gate_1582(n1610,n1606,n1609);
not gate_1583(n1611,n1610);
and gate_1584(n1612,pi7,n1611);
not gate_1585(n1613,n1612);
and gate_1586(n1614,n31,n1182);
and gate_1587(n1615,n129,n1614);
not gate_1588(n1616,n1615);
and gate_1589(n1617,n1613,n1616);
not gate_1590(n1618,n1617);
and gate_1591(n1619,pi0,n1618);
not gate_1592(n1620,n1619);
and gate_1593(n1621,n1600,n1620);
and gate_1594(n1622,n1526,n1621);
not gate_1595(n1623,n1622);
and gate_1596(n1624,n36,n1623);
not gate_1597(n1625,n1624);
and gate_1598(n1626,pi1,n1188);
not gate_1599(n1627,n1626);
and gate_1600(n1628,n299,n662);
not gate_1601(n1629,n1628);
and gate_1602(n1630,n1627,n1629);
not gate_1603(n1631,n1630);
and gate_1604(n1632,n35,n1631);
not gate_1605(n1633,n1632);
and gate_1606(n1634,pi4,n590);
not gate_1607(n1635,n1634);
and gate_1608(n1636,n1241,n1634);
not gate_1609(n1637,n1636);
and gate_1610(n1638,n1633,n1637);
not gate_1611(n1639,n1638);
and gate_1612(n1640,pi3,n1639);
not gate_1613(n1641,n1640);
and gate_1614(n1642,pi1,n1154);
and gate_1615(n1643,n811,n1642);
not gate_1616(n1644,n1643);
and gate_1617(n1645,n1641,n1644);
not gate_1618(n1646,n1645);
and gate_1619(n1647,pi7,n1646);
not gate_1620(n1648,n1647);
and gate_1621(n1649,n32,n662);
not gate_1622(n1650,n1649);
and gate_1623(n1651,n1508,n1650);
not gate_1624(n1652,n1651);
and gate_1625(n1653,pi5,n1652);
and gate_1626(n1654,pi1,n202);
and gate_1627(n1655,n1653,n1654);
not gate_1628(n1656,n1655);
and gate_1629(n1657,n1648,n1656);
not gate_1630(n1658,n1657);
and gate_1631(n1659,pi0,n1658);
not gate_1632(n1660,n1659);
and gate_1633(n1661,n1625,n1660);
and gate_1634(n1662,n1449,n1661);
and gate_1635(n1663,n1268,n1662);
not gate_1636(po04,n1663);
and gate_1637(n1665,pi0,n1145);
and gate_1638(n1666,n206,n1078);
and gate_1639(n1667,n1665,n1666);
not gate_1640(n1668,n1667);
and gate_1641(n1669,n706,n1259);
not gate_1642(n1670,n1669);
and gate_1643(n1671,pi0,n1131);
and gate_1644(n1672,n34,n1671);
not gate_1645(n1673,n1672);
and gate_1646(n1674,n1670,n1673);
not gate_1647(n1675,n1674);
and gate_1648(n1676,pi3,n1675);
not gate_1649(n1677,n1676);
and gate_1650(n1678,n1668,n1677);
not gate_1651(n1679,n1678);
and gate_1652(n1680,n421,n1679);
not gate_1653(n1681,n1680);
and gate_1654(n1682,n597,n1635);
not gate_1655(n1683,n1682);
and gate_1656(n1684,pi0,n1683);
not gate_1657(n1685,n1684);
and gate_1658(n1686,n455,n768);
not gate_1659(n1687,n1686);
and gate_1660(n1688,n1685,n1687);
not gate_1661(n1689,n1688);
and gate_1662(n1690,pi3,n1689);
not gate_1663(n1691,n1690);
and gate_1664(n1692,n30,n33);
not gate_1665(n1693,n1692);
and gate_1666(n1694,n572,n1692);
not gate_1667(n1695,n1694);
and gate_1668(n1696,n1691,n1695);
not gate_1669(n1697,n1696);
and gate_1670(n1698,pi1,n1697);
not gate_1671(n1699,n1698);
and gate_1672(n1700,pi0,n980);
not gate_1673(n1701,n1700);
and gate_1674(n1702,n143,n164);
and gate_1675(n1703,n637,n1702);
and gate_1676(n1704,n1700,n1703);
not gate_1677(n1705,n1704);
and gate_1678(n1706,n1699,n1705);
not gate_1679(n1707,n1706);
and gate_1680(n1708,n32,n1707);
not gate_1681(n1709,n1708);
and gate_1682(n1710,pi0,pi3);
and gate_1683(n1711,n1634,n1710);
not gate_1684(n1712,n1711);
and gate_1685(n1713,n816,n1692);
not gate_1686(n1714,n1713);
and gate_1687(n1715,n1712,n1714);
not gate_1688(n1716,n1715);
and gate_1689(n1717,n31,n1716);
not gate_1690(n1718,n1717);
and gate_1691(n1719,n1494,n1710);
not gate_1692(n1720,n1719);
and gate_1693(n1721,n1718,n1720);
not gate_1694(n1722,n1721);
and gate_1695(n1723,pi2,n1722);
not gate_1696(n1724,n1723);
and gate_1697(n1725,n1709,n1724);
not gate_1698(n1726,n1725);
and gate_1699(n1727,pi6,n1726);
not gate_1700(n1728,n1727);
and gate_1701(n1729,n817,n1586);
not gate_1702(n1730,n1729);
and gate_1703(n1731,n277,n336);
not gate_1704(n1732,n1731);
and gate_1705(n1733,n1729,n1731);
not gate_1706(n1734,n1733);
and gate_1707(n1735,n1728,n1734);
and gate_1708(n1736,pi4,n1007);
not gate_1709(n1737,n1736);
and gate_1710(n1738,n34,n1078);
not gate_1711(n1739,n1738);
and gate_1712(n1740,n1737,n1739);
not gate_1713(n1741,n1740);
and gate_1714(n1742,n140,n1741);
not gate_1715(n1743,n1742);
and gate_1716(n1744,n427,n694);
and gate_1717(n1745,n30,n1744);
not gate_1718(n1746,n1745);
and gate_1719(n1747,n1743,n1746);
not gate_1720(n1748,n1747);
and gate_1721(n1749,n38,n1748);
not gate_1722(n1750,n1749);
and gate_1723(n1751,n97,n285);
not gate_1724(n1752,n1751);
and gate_1725(n1753,pi6,n707);
and gate_1726(n1754,pi4,n1004);
not gate_1727(n1755,n1754);
and gate_1728(n1756,n1753,n1755);
not gate_1729(n1757,n1756);
and gate_1730(n1758,n1752,n1757);
not gate_1731(n1759,n1758);
and gate_1732(n1760,n30,n1759);
not gate_1733(n1761,n1760);
and gate_1734(n1762,pi0,n34);
and gate_1735(n1763,n106,n1762);
not gate_1736(n1764,n1763);
and gate_1737(n1765,n1761,n1764);
not gate_1738(n1766,n1765);
and gate_1739(n1767,pi8,n1766);
not gate_1740(n1768,n1767);
and gate_1741(n1769,n1750,n1768);
not gate_1742(n1770,n1769);
and gate_1743(n1771,pi1,n1770);
not gate_1744(n1772,n1771);
and gate_1745(n1773,n250,n456);
not gate_1746(n1774,n1773);
and gate_1747(n1775,pi7,n1774);
not gate_1748(n1776,n1775);
and gate_1749(n1777,n130,n1776);
not gate_1750(n1778,n1777);
and gate_1751(n1779,n36,n1778);
not gate_1752(n1780,n1779);
and gate_1753(n1781,pi7,n1195);
not gate_1754(n1782,n1781);
and gate_1755(n1783,n150,n1782);
not gate_1756(n1784,n1783);
and gate_1757(n1785,n1780,n1784);
not gate_1758(n1786,n1785);
and gate_1759(n1787,pi0,n1786);
not gate_1760(n1788,n1787);
and gate_1761(n1789,pi8,n1128);
and gate_1762(n1790,n1155,n1789);
not gate_1763(n1791,n1790);
and gate_1764(n1792,n1788,n1791);
not gate_1765(n1793,n1792);
and gate_1766(n1794,n34,n1793);
not gate_1767(n1795,n1794);
and gate_1768(n1796,n39,n137);
not gate_1769(n1797,n1796);
and gate_1770(n1798,n35,n88);
not gate_1771(n1799,n1798);
and gate_1772(n1800,pi7,n1799);
not gate_1773(n1801,n1800);
and gate_1774(n1802,n999,n1801);
not gate_1775(n1803,n1802);
and gate_1776(n1804,n38,n1803);
not gate_1777(n1805,n1804);
and gate_1778(n1806,n39,n150);
not gate_1779(n1807,n1806);
and gate_1780(n1808,n1805,n1807);
not gate_1781(n1809,n1808);
and gate_1782(n1810,n768,n1809);
not gate_1783(n1811,n1810);
and gate_1784(n1812,n1797,n1811);
not gate_1785(n1813,n1812);
and gate_1786(n1814,n31,n1813);
not gate_1787(n1815,n1814);
and gate_1788(n1816,n1795,n1815);
and gate_1789(n1817,n1772,n1816);
not gate_1790(n1818,n1817);
and gate_1791(n1819,pi3,n1818);
not gate_1792(n1820,n1819);
and gate_1793(n1821,n81,n175);
not gate_1794(n1822,n1821);
and gate_1795(n1823,n53,n87);
not gate_1796(n1824,n1823);
and gate_1797(n1825,n1822,n1824);
not gate_1798(n1826,n1825);
and gate_1799(n1827,pi0,n1826);
not gate_1800(n1828,n1827);
and gate_1801(n1829,n30,pi5);
and gate_1802(n1830,n54,n333);
not gate_1803(n1831,n1830);
and gate_1804(n1832,n1829,n1831);
not gate_1805(n1833,n1832);
and gate_1806(n1834,n149,n1833);
and gate_1807(n1835,n1828,n1834);
not gate_1808(n1836,n1835);
and gate_1809(n1837,pi4,n1836);
not gate_1810(n1838,n1837);
and gate_1811(n1839,pi0,n919);
not gate_1812(n1840,n1839);
and gate_1813(n1841,pi0,n37);
not gate_1814(n1842,n1841);
and gate_1815(n1843,n190,n1842);
and gate_1816(n1844,n636,n1843);
not gate_1817(n1845,n1844);
and gate_1818(n1846,n1840,n1845);
not gate_1819(n1847,n1846);
and gate_1820(n1848,pi5,n1847);
not gate_1821(n1849,n1848);
and gate_1822(n1850,n40,n958);
not gate_1823(n1851,n1850);
and gate_1824(n1852,n30,n1851);
not gate_1825(n1853,n1852);
and gate_1826(n1854,n35,n53);
not gate_1827(n1855,n1854);
and gate_1828(n1856,n1853,n1855);
not gate_1829(n1857,n1856);
and gate_1830(n1858,n784,n1857);
not gate_1831(n1859,n1858);
and gate_1832(n1860,n1849,n1859);
and gate_1833(n1861,n1838,n1860);
not gate_1834(n1862,n1861);
and gate_1835(n1863,pi1,n1862);
not gate_1836(n1864,n1863);
and gate_1837(n1865,n332,n608);
not gate_1838(n1866,n1865);
and gate_1839(n1867,n176,n1866);
not gate_1840(n1868,n1867);
and gate_1841(n1869,n37,n1868);
not gate_1842(n1870,n1869);
and gate_1843(n1871,pi5,n336);
not gate_1844(n1872,n1871);
and gate_1845(n1873,n729,n1872);
not gate_1846(n1874,n1873);
and gate_1847(n1875,pi4,n1874);
not gate_1848(n1876,n1875);
and gate_1849(n1877,n35,n336);
not gate_1850(n1878,n1877);
and gate_1851(n1879,n151,n1878);
not gate_1852(n1880,n1879);
and gate_1853(n1881,n34,n1880);
not gate_1854(n1882,n1881);
and gate_1855(n1883,n1876,n1882);
not gate_1856(n1884,n1883);
and gate_1857(n1885,pi7,n1884);
not gate_1858(n1886,n1885);
and gate_1859(n1887,n285,n358);
not gate_1860(n1888,n1887);
and gate_1861(n1889,n1886,n1888);
and gate_1862(n1890,n1870,n1889);
not gate_1863(n1891,n1890);
and gate_1864(n1892,pi0,n1891);
not gate_1865(n1893,n1892);
and gate_1866(n1894,n39,n277);
not gate_1867(n1895,n1894);
and gate_1868(n1896,n135,n1894);
not gate_1869(n1897,n1896);
and gate_1870(n1898,n1893,n1897);
not gate_1871(n1899,n1898);
and gate_1872(n1900,n31,n1899);
not gate_1873(n1901,n1900);
and gate_1874(n1902,n1864,n1901);
not gate_1875(n1903,n1902);
and gate_1876(n1904,n33,n1903);
not gate_1877(n1905,n1904);
and gate_1878(n1906,n66,n838);
not gate_1879(n1907,n1906);
and gate_1880(n1908,n31,n509);
not gate_1881(n1909,n1908);
and gate_1882(n1910,n1907,n1908);
and gate_1883(n1911,pi0,n1910);
not gate_1884(n1912,n1911);
and gate_1885(n1913,n1905,n1912);
and gate_1886(n1914,n1820,n1913);
not gate_1887(n1915,n1914);
and gate_1888(n1916,pi2,n1915);
not gate_1889(n1917,n1916);
and gate_1890(n1918,n32,n36);
not gate_1891(n1919,n1918);
and gate_1892(n1920,n115,n1918);
not gate_1893(n1921,n1920);
and gate_1894(n1922,n226,n1921);
not gate_1895(n1923,n1922);
and gate_1896(n1924,n37,n1923);
not gate_1897(n1925,n1924);
and gate_1898(n1926,n32,n146);
not gate_1899(n1927,n1926);
and gate_1900(n1928,n997,n1927);
not gate_1901(n1929,n1928);
and gate_1902(n1930,n33,n1929);
not gate_1903(n1931,n1930);
and gate_1904(n1932,n1925,n1931);
not gate_1905(n1933,n1932);
and gate_1906(n1934,n38,n1933);
not gate_1907(n1935,n1934);
and gate_1908(n1936,n33,n39);
not gate_1909(n1937,n1936);
and gate_1910(n1938,pi2,n147);
not gate_1911(n1939,n1938);
and gate_1912(n1940,n1936,n1939);
not gate_1913(n1941,n1940);
and gate_1914(n1942,n1935,n1941);
not gate_1915(n1943,n1942);
and gate_1916(n1944,n34,n1943);
not gate_1917(n1945,n1944);
and gate_1918(n1946,n181,n218);
not gate_1919(n1947,n1946);
and gate_1920(n1948,n179,n240);
not gate_1921(n1949,n1948);
and gate_1922(n1950,n1947,n1949);
not gate_1923(n1951,n1950);
and gate_1924(n1952,pi8,n1951);
not gate_1925(n1953,n1952);
and gate_1926(n1954,pi3,n175);
not gate_1927(n1955,n1954);
and gate_1928(n1956,n90,n1955);
not gate_1929(n1957,n1956);
and gate_1930(n1958,n43,n1957);
not gate_1931(n1959,n1958);
and gate_1932(n1960,n1953,n1959);
not gate_1933(n1961,n1960);
and gate_1934(n1962,n32,n1961);
not gate_1935(n1963,n1962);
and gate_1936(n1964,n217,n617);
not gate_1937(n1965,n1964);
and gate_1938(n1966,n1963,n1965);
not gate_1939(n1967,n1966);
and gate_1940(n1968,pi4,n1967);
not gate_1941(n1969,n1968);
and gate_1942(n1970,n1945,n1969);
not gate_1943(n1971,n1970);
and gate_1944(n1972,n31,n1971);
not gate_1945(n1973,n1972);
and gate_1946(n1974,n258,n1325);
not gate_1947(n1975,n1974);
and gate_1948(n1976,pi3,n1975);
not gate_1949(n1977,n1976);
and gate_1950(n1978,n33,n884);
not gate_1951(n1979,n1978);
and gate_1952(n1980,n1977,n1979);
not gate_1953(n1981,n1980);
and gate_1954(n1982,n36,n1981);
not gate_1955(n1983,n1982);
and gate_1956(n1984,n51,n885);
not gate_1957(n1985,n1984);
and gate_1958(n1986,n1983,n1985);
not gate_1959(n1987,n1986);
and gate_1960(n1988,n38,n1987);
not gate_1961(n1989,n1988);
and gate_1962(n1990,n310,n627);
not gate_1963(n1991,n1990);
and gate_1964(n1992,n81,n1991);
not gate_1965(n1993,n1992);
and gate_1966(n1994,n1989,n1993);
not gate_1967(n1995,n1994);
and gate_1968(n1996,pi5,n1995);
not gate_1969(n1997,n1996);
and gate_1970(n1998,n310,n631);
and gate_1971(n1999,n906,n1998);
not gate_1972(n2000,n1999);
and gate_1973(n2001,pi4,n2000);
not gate_1974(n2002,n2001);
and gate_1975(n2003,n142,n666);
not gate_1976(n2004,n2003);
and gate_1977(n2005,n2002,n2004);
not gate_1978(n2006,n2005);
and gate_1979(n2007,n35,n2006);
not gate_1980(n2008,n2007);
and gate_1981(n2009,n1997,n2008);
not gate_1982(n2010,n2009);
and gate_1983(n2011,pi1,n2010);
not gate_1984(n2012,n2011);
and gate_1985(n2013,n41,n465);
not gate_1986(n2014,n2013);
and gate_1987(n2015,n2012,n2014);
not gate_1988(n2016,n2015);
and gate_1989(n2017,n32,n2016);
not gate_1990(n2018,n2017);
and gate_1991(n2019,n1973,n2018);
not gate_1992(n2020,n2019);
and gate_1993(n2021,pi0,n2020);
not gate_1994(n2022,n2021);
and gate_1995(n2023,pi4,n87);
not gate_1996(n2024,n2023);
and gate_1997(n2025,n510,n2024);
not gate_1998(n2026,n2025);
and gate_1999(n2027,n260,n2026);
not gate_2000(n2028,n2027);
and gate_2001(n2029,n104,n277);
not gate_2002(n2030,n2029);
and gate_2003(n2031,n999,n2030);
not gate_2004(n2032,n2031);
and gate_2005(n2033,pi8,n2032);
not gate_2006(n2034,n2033);
and gate_2007(n2035,n2028,n2034);
not gate_2008(n2036,n2035);
and gate_2009(n2037,n33,n2036);
not gate_2010(n2038,n2037);
and gate_2011(n2039,n34,n150);
not gate_2012(n2040,n2039);
and gate_2013(n2041,n745,n2040);
not gate_2014(n2042,n2041);
and gate_2015(n2043,pi8,n178);
and gate_2016(n2044,pi4,n2043);
not gate_2017(n2045,n2044);
and gate_2018(n2046,n2041,n2045);
not gate_2019(n2047,n2046);
and gate_2020(n2048,n37,n2047);
not gate_2021(n2049,n2048);
and gate_2022(n2050,pi8,n419);
not gate_2023(n2051,n2050);
and gate_2024(n2052,n34,n2051);
not gate_2025(n2053,n2052);
and gate_2026(n2054,n337,n2053);
not gate_2027(n2055,n2054);
and gate_2028(n2056,pi7,n2055);
not gate_2029(n2057,n2056);
and gate_2030(n2058,n82,n626);
not gate_2031(n2059,n2058);
and gate_2032(n2060,n2057,n2059);
not gate_2033(n2061,n2060);
and gate_2034(n2062,n35,n2061);
not gate_2035(n2063,n2062);
and gate_2036(n2064,n104,n509);
not gate_2037(n2065,n2064);
and gate_2038(n2066,n2063,n2065);
and gate_2039(n2067,n2049,n2066);
not gate_2040(n2068,n2067);
and gate_2041(n2069,pi3,n2068);
not gate_2042(n2070,n2069);
and gate_2043(n2071,n2038,n2070);
not gate_2044(n2072,n2071);
and gate_2045(n2073,n32,n2072);
not gate_2046(n2074,n2073);
and gate_2047(n2075,n65,n542);
not gate_2048(n2076,n2075);
and gate_2049(n2077,n2074,n2076);
not gate_2050(n2078,n2077);
and gate_2051(n2079,n30,n2078);
not gate_2052(n2080,n2079);
and gate_2053(n2081,n32,n206);
and gate_2054(n2082,n724,n2081);
not gate_2055(n2083,n2082);
and gate_2056(n2084,n2080,n2083);
not gate_2057(n2085,n2084);
and gate_2058(n2086,pi1,n2085);
not gate_2059(n2087,n2086);
and gate_2060(n2088,n2022,n2087);
and gate_2061(n2089,n1917,n2088);
and gate_2062(n2090,n1735,n2089);
and gate_2063(n2091,n1681,n2090);
not gate_2064(po05,n2091);
and gate_2065(n2093,pi0,n32);
and gate_2066(n2094,n192,n2093);
not gate_2067(n2095,n2094);
and gate_2068(n2096,n1320,n2095);
not gate_2069(n2097,n2096);
and gate_2070(n2098,n35,n2097);
not gate_2071(n2099,n2098);
and gate_2072(n2100,pi3,n509);
and gate_2073(n2101,n2093,n2100);
not gate_2074(n2102,n2101);
and gate_2075(n2103,n2099,n2102);
not gate_2076(n2104,n2103);
and gate_2077(n2105,pi6,n2104);
not gate_2078(n2106,n2105);
and gate_2079(n2107,n1215,n1954);
not gate_2080(n2108,n2107);
and gate_2081(n2109,n2106,n2108);
not gate_2082(n2110,n2109);
and gate_2083(n2111,pi1,n2110);
not gate_2084(n2112,n2111);
and gate_2085(n2113,n34,n87);
and gate_2086(n2114,n69,n2113);
not gate_2087(n2115,n2114);
and gate_2088(n2116,n768,n1954);
not gate_2089(n2117,n2116);
and gate_2090(n2118,n2115,n2117);
not gate_2091(n2119,n2118);
and gate_2092(n2120,pi2,n2119);
not gate_2093(n2121,n2120);
and gate_2094(n2122,n33,n626);
not gate_2095(n2123,n2122);
and gate_2096(n2124,n2093,n2122);
not gate_2097(n2125,n2124);
and gate_2098(n2126,n2121,n2125);
not gate_2099(n2127,n2126);
and gate_2100(n2128,n31,n2127);
not gate_2101(n2129,n2128);
and gate_2102(n2130,n2112,n2129);
not gate_2103(n2131,n2130);
and gate_2104(n2132,pi8,n2131);
not gate_2105(n2133,n2132);
and gate_2106(n2134,n1138,n1242);
not gate_2107(n2135,n2134);
and gate_2108(n2136,n2023,n2135);
and gate_2109(n2137,pi0,n2136);
not gate_2110(n2138,n2137);
and gate_2111(n2139,n34,n175);
and gate_2112(n2140,n1259,n2139);
not gate_2113(n2141,n2140);
and gate_2114(n2142,n2138,n2141);
not gate_2115(n2143,n2142);
and gate_2116(n2144,pi3,n2143);
not gate_2117(n2145,n2144);
and gate_2118(n2146,n30,n87);
not gate_2119(n2147,n2146);
and gate_2120(n2148,n206,n299);
not gate_2121(n2149,n2148);
and gate_2122(n2150,n2146,n2148);
not gate_2123(n2151,n2150);
and gate_2124(n2152,n2145,n2151);
not gate_2125(n2153,n2152);
and gate_2126(n2154,n38,n2153);
not gate_2127(n2155,n2154);
and gate_2128(n2156,n2133,n2155);
and gate_2129(n2157,n151,n529);
not gate_2130(n2158,n2157);
and gate_2131(n2159,pi4,n2158);
not gate_2132(n2160,n2159);
and gate_2133(n2161,n454,n456);
not gate_2134(n2162,n2161);
and gate_2135(n2163,n424,n2162);
not gate_2136(n2164,n2163);
and gate_2137(n2165,n1872,n2164);
and gate_2138(n2166,n2160,n2165);
not gate_2139(n2167,n2166);
and gate_2140(n2168,pi1,n2167);
not gate_2141(n2169,n2168);
and gate_2142(n2170,n285,n332);
not gate_2143(n2171,n2170);
and gate_2144(n2172,n35,n785);
not gate_2145(n2173,n2172);
and gate_2146(n2174,pi5,n784);
not gate_2147(n2175,n2174);
and gate_2148(n2176,n2173,n2175);
and gate_2149(n2177,n38,n2176);
not gate_2150(n2178,n2177);
and gate_2151(n2179,n2171,n2178);
not gate_2152(n2180,n2179);
and gate_2153(n2181,n31,n2180);
not gate_2154(n2182,n2181);
and gate_2155(n2183,n2169,n2182);
not gate_2156(n2184,n2183);
and gate_2157(n2185,n30,n2184);
not gate_2158(n2186,n2185);
and gate_2159(n2187,n31,n1156);
not gate_2160(n2188,n2187);
and gate_2161(n2189,pi8,n2188);
not gate_2162(n2190,n2189);
and gate_2163(n2191,n31,n358);
not gate_2164(n2192,n2191);
and gate_2165(n2193,n2190,n2192);
not gate_2166(n2194,n2193);
and gate_2167(n2195,pi5,n2194);
not gate_2168(n2196,n2195);
and gate_2169(n2197,n333,n337);
not gate_2170(n2198,n2197);
and gate_2171(n2199,pi1,n2198);
not gate_2172(n2200,n2199);
and gate_2173(n2201,n419,n2200);
not gate_2174(n2202,n2201);
and gate_2175(n2203,n35,n2202);
not gate_2176(n2204,n2203);
and gate_2177(n2205,n2196,n2204);
not gate_2178(n2206,n2205);
and gate_2179(n2207,n34,n2206);
not gate_2180(n2208,n2207);
and gate_2181(n2209,n31,n422);
not gate_2182(n2210,n2209);
and gate_2183(n2211,pi1,n358);
not gate_2184(n2212,n2211);
and gate_2185(n2213,n2210,n2212);
not gate_2186(n2214,n2213);
and gate_2187(n2215,pi5,n2214);
not gate_2188(n2216,n2215);
and gate_2189(n2217,n2208,n2216);
not gate_2190(n2218,n2217);
and gate_2191(n2219,pi0,n2218);
not gate_2192(n2220,n2219);
and gate_2193(n2221,n2186,n2220);
not gate_2194(n2222,n2221);
and gate_2195(n2223,pi3,n2222);
not gate_2196(n2224,n2223);
and gate_2197(n2225,n313,n332);
not gate_2198(n2226,n2225);
and gate_2199(n2227,n139,n419);
not gate_2200(n2228,n2227);
and gate_2201(n2229,pi1,n2228);
not gate_2202(n2230,n2229);
and gate_2203(n2231,n2226,n2230);
not gate_2204(n2232,n2231);
and gate_2205(n2233,n34,n2232);
not gate_2206(n2234,n2233);
and gate_2207(n2235,pi0,n2191);
not gate_2208(n2236,n2235);
and gate_2209(n2237,n314,n418);
not gate_2210(n2238,n2237);
and gate_2211(n2239,n2236,n2238);
not gate_2212(n2240,n2239);
and gate_2213(n2241,pi4,n2240);
not gate_2214(n2242,n2241);
and gate_2215(n2243,pi0,n31);
not gate_2216(n2244,n2243);
and gate_2217(n2245,n336,n2243);
not gate_2218(n2246,n2245);
and gate_2219(n2247,n2242,n2246);
and gate_2220(n2248,n2234,n2247);
not gate_2221(n2249,n2248);
and gate_2222(n2250,pi5,n2249);
not gate_2223(n2251,n2250);
and gate_2224(n2252,n347,n627);
not gate_2225(n2253,n2252);
and gate_2226(n2254,n769,n2253);
and gate_2227(n2255,pi1,n2254);
not gate_2228(n2256,n2255);
and gate_2229(n2257,pi4,n336);
not gate_2230(n2258,n2257);
and gate_2231(n2259,n2243,n2257);
not gate_2232(n2260,n2259);
and gate_2233(n2261,n2256,n2260);
not gate_2234(n2262,n2261);
and gate_2235(n2263,n35,n2262);
not gate_2236(n2264,n2263);
and gate_2237(n2265,n2251,n2264);
not gate_2238(n2266,n2265);
and gate_2239(n2267,n33,n2266);
not gate_2240(n2268,n2267);
and gate_2241(n2269,n423,n453);
and gate_2242(n2270,n2243,n2269);
not gate_2243(n2271,n2270);
and gate_2244(n2272,n2268,n2271);
and gate_2245(n2273,n2224,n2272);
not gate_2246(n2274,n2273);
and gate_2247(n2275,n37,n2274);
not gate_2248(n2276,n2275);
and gate_2249(n2277,n522,n2258);
not gate_2250(n2278,n2277);
and gate_2251(n2279,n207,n2278);
and gate_2252(n2280,pi0,n2279);
not gate_2253(n2281,n2280);
and gate_2254(n2282,n385,n768);
not gate_2255(n2283,n2282);
and gate_2256(n2284,n2281,n2283);
and gate_2257(n2285,pi5,n332);
not gate_2258(n2286,n2285);
and gate_2259(n2287,n785,n2286);
not gate_2260(n2288,n2287);
and gate_2261(n2289,n33,n2288);
not gate_2262(n2290,n2289);
and gate_2263(n2291,pi5,n591);
not gate_2264(n2292,n2291);
and gate_2265(n2293,n424,n2292);
and gate_2266(n2294,pi3,n2293);
not gate_2267(n2295,n2294);
and gate_2268(n2296,n52,n177);
and gate_2269(n2297,n451,n2296);
not gate_2270(n2298,n2297);
and gate_2271(n2299,n2295,n2298);
and gate_2272(n2300,n2290,n2299);
not gate_2273(n2301,n2300);
and gate_2274(n2302,n30,n2301);
not gate_2275(n2303,n2302);
and gate_2276(n2304,pi4,n150);
not gate_2277(n2305,n2304);
and gate_2278(n2306,n573,n2305);
not gate_2279(n2307,n2306);
and gate_2280(n2308,pi3,n2307);
not gate_2281(n2309,n2308);
and gate_2282(n2310,n206,n358);
not gate_2283(n2311,n2310);
and gate_2284(n2312,n2309,n2311);
not gate_2285(n2313,n2312);
and gate_2286(n2314,pi0,n2313);
not gate_2287(n2315,n2314);
and gate_2288(n2316,n2303,n2315);
and gate_2289(n2317,n2284,n2316);
not gate_2290(n2318,n2317);
and gate_2291(n2319,pi1,n2318);
not gate_2292(n2320,n2319);
and gate_2293(n2321,n418,n768);
not gate_2294(n2322,n2321);
and gate_2295(n2323,pi0,pi4);
not gate_2296(n2324,n2323);
and gate_2297(n2325,n1553,n2324);
not gate_2298(n2326,n2325);
and gate_2299(n2327,n38,n2325);
and gate_2300(n2328,n423,n2327);
not gate_2301(n2329,n2328);
and gate_2302(n2330,n2322,n2329);
not gate_2303(n2331,n2330);
and gate_2304(n2332,n35,n2331);
not gate_2305(n2333,n2332);
and gate_2306(n2334,n30,n332);
not gate_2307(n2335,n2334);
and gate_2308(n2336,n336,n2323);
not gate_2309(n2337,n2336);
and gate_2310(n2338,n2335,n2337);
not gate_2311(n2339,n2338);
and gate_2312(n2340,pi5,n2339);
not gate_2313(n2341,n2340);
and gate_2314(n2342,n2333,n2341);
not gate_2315(n2343,n2342);
and gate_2316(n2344,pi3,n2343);
not gate_2317(n2345,n2344);
and gate_2318(n2346,n69,n99);
not gate_2319(n2347,n2346);
and gate_2320(n2348,n30,n590);
not gate_2321(n2349,n2348);
and gate_2322(n2350,n2347,n2349);
not gate_2323(n2351,n2350);
and gate_2324(n2352,pi4,n2351);
not gate_2325(n2353,n2352);
and gate_2326(n2354,n510,n749);
not gate_2327(n2355,n2354);
and gate_2328(n2356,n345,n2355);
and gate_2329(n2357,pi0,n2356);
not gate_2330(n2358,n2357);
and gate_2331(n2359,n2353,n2358);
not gate_2332(n2360,n2359);
and gate_2333(n2361,pi6,n2360);
not gate_2334(n2362,n2361);
and gate_2335(n2363,pi0,n142);
and gate_2336(n2364,n1877,n2363);
not gate_2337(n2365,n2364);
and gate_2338(n2366,n2362,n2365);
and gate_2339(n2367,n2345,n2366);
not gate_2340(n2368,n2367);
and gate_2341(n2369,n31,n2368);
not gate_2342(n2370,n2369);
and gate_2343(n2371,n777,n1216);
not gate_2344(n2372,n2371);
and gate_2345(n2373,n2370,n2372);
and gate_2346(n2374,n2320,n2373);
not gate_2347(n2375,n2374);
and gate_2348(n2376,pi7,n2375);
not gate_2349(n2377,n2376);
and gate_2350(n2378,n636,n1710);
not gate_2351(n2379,n2378);
and gate_2352(n2380,n33,n455);
and gate_2353(n2381,n768,n2380);
not gate_2354(n2382,n2381);
and gate_2355(n2383,n2379,n2382);
not gate_2356(n2384,n2383);
and gate_2357(n2385,pi6,n2384);
and gate_2358(n2386,pi1,n2385);
not gate_2359(n2387,n2386);
and gate_2360(n2388,n2377,n2387);
and gate_2361(n2389,n2276,n2388);
not gate_2362(n2390,n2389);
and gate_2363(n2391,pi2,n2390);
not gate_2364(n2392,n2391);
and gate_2365(n2393,n1732,n1866);
not gate_2366(n2394,n2393);
and gate_2367(n2395,pi0,pi1);
not gate_2368(n2396,n2395);
and gate_2369(n2397,n314,n2396);
not gate_2370(n2398,n2397);
and gate_2371(n2399,n31,n219);
not gate_2372(n2400,n2399);
and gate_2373(n2401,n222,n2400);
not gate_2374(n2402,n2401);
and gate_2375(n2403,n2397,n2402);
and gate_2376(n2404,n2394,n2403);
not gate_2377(n2405,n2404);
and gate_2378(n2406,n163,n728);
not gate_2379(n2407,n2406);
and gate_2380(n2408,n336,n509);
not gate_2381(n2409,n2408);
and gate_2382(n2410,n2407,n2409);
not gate_2383(n2411,n2410);
and gate_2384(n2412,n31,n2411);
not gate_2385(n2413,n2412);
and gate_2386(n2414,n609,n1217);
and gate_2387(n2415,n278,n358);
not gate_2388(n2416,n2415);
and gate_2389(n2417,n2414,n2416);
and gate_2390(n2418,n33,n2417);
not gate_2391(n2419,n2418);
and gate_2392(n2420,n456,n595);
not gate_2393(n2421,n2420);
and gate_2394(n2422,n36,n2421);
not gate_2395(n2423,n2422);
and gate_2396(n2424,n358,n608);
not gate_2397(n2425,n2424);
and gate_2398(n2426,n2423,n2425);
not gate_2399(n2427,n2426);
and gate_2400(n2428,pi3,n2427);
not gate_2401(n2429,n2428);
and gate_2402(n2430,n2419,n2429);
not gate_2403(n2431,n2430);
and gate_2404(n2432,pi1,n2431);
not gate_2405(n2433,n2432);
and gate_2406(n2434,n163,n1216);
not gate_2407(n2435,n2434);
and gate_2408(n2436,n142,n931);
not gate_2409(n2437,n2436);
and gate_2410(n2438,n2435,n2437);
and gate_2411(n2439,n2433,n2438);
and gate_2412(n2440,n2413,n2439);
not gate_2413(n2441,n2440);
and gate_2414(n2442,pi7,n2441);
not gate_2415(n2443,n2442);
and gate_2416(n2444,n435,n455);
not gate_2417(n2445,n2444);
and gate_2418(n2446,n1495,n2445);
not gate_2419(n2447,n2446);
and gate_2420(n2448,n312,n2447);
not gate_2421(n2449,n2448);
and gate_2422(n2450,n1253,n1355);
and gate_2423(n2451,n143,n2450);
and gate_2424(n2452,pi1,n2451);
not gate_2425(n2453,n2452);
and gate_2426(n2454,n749,n812);
not gate_2427(n2455,n2454);
and gate_2428(n2456,n207,n2455);
and gate_2429(n2457,n31,n2456);
not gate_2430(n2458,n2457);
and gate_2431(n2459,n142,n453);
not gate_2432(n2460,n2459);
and gate_2433(n2461,n2458,n2460);
and gate_2434(n2462,n2453,n2461);
not gate_2435(n2463,n2462);
and gate_2436(n2464,n36,n2463);
not gate_2437(n2465,n2464);
and gate_2438(n2466,n590,n799);
not gate_2439(n2467,n2466);
and gate_2440(n2468,n520,n1534);
not gate_2441(n2469,n2468);
and gate_2442(n2470,n2467,n2469);
not gate_2443(n2471,n2470);
and gate_2444(n2472,n626,n2471);
not gate_2445(n2473,n2472);
and gate_2446(n2474,n2465,n2473);
and gate_2447(n2475,n2449,n2474);
not gate_2448(n2476,n2475);
and gate_2449(n2477,n37,n2476);
not gate_2450(n2478,n2477);
and gate_2451(n2479,n31,n142);
and gate_2452(n2480,n1877,n2479);
not gate_2453(n2481,n2480);
and gate_2454(n2482,n2478,n2481);
and gate_2455(n2483,n2443,n2482);
not gate_2456(n2484,n2483);
and gate_2457(n2485,pi0,n2484);
not gate_2458(n2486,n2485);
and gate_2459(n2487,n34,n358);
not gate_2460(n2488,n2487);
and gate_2461(n2489,n529,n2488);
not gate_2462(n2490,n2489);
and gate_2463(n2491,n609,n2490);
and gate_2464(n2492,n33,n2491);
not gate_2465(n2493,n2492);
and gate_2466(n2494,n583,n2198);
not gate_2467(n2495,n2494);
and gate_2468(n2496,n150,n639);
not gate_2469(n2497,n2496);
and gate_2470(n2498,n2495,n2497);
not gate_2471(n2499,n2498);
and gate_2472(n2500,pi3,n2499);
not gate_2473(n2501,n2500);
and gate_2474(n2502,n2493,n2501);
not gate_2475(n2503,n2502);
and gate_2476(n2504,n37,n2503);
not gate_2477(n2505,n2504);
and gate_2478(n2506,n418,n509);
not gate_2479(n2507,n2506);
and gate_2480(n2508,n2024,n2507);
not gate_2481(n2509,n2508);
and gate_2482(n2510,pi7,n2509);
not gate_2483(n2511,n2510);
and gate_2484(n2512,n2409,n2511);
not gate_2485(n2513,n2512);
and gate_2486(n2514,n33,n2513);
not gate_2487(n2515,n2514);
and gate_2488(n2516,n35,n179);
not gate_2489(n2517,n2516);
and gate_2490(n2518,pi4,n1753);
not gate_2491(n2519,n2518);
and gate_2492(n2520,n2517,n2519);
not gate_2493(n2521,n2520);
and gate_2494(n2522,n38,n2521);
not gate_2495(n2523,n2522);
and gate_2496(n2524,n418,n608);
not gate_2497(n2525,n2524);
and gate_2498(n2526,n2523,n2525);
not gate_2499(n2527,n2526);
and gate_2500(n2528,pi3,n2527);
not gate_2501(n2529,n2528);
and gate_2502(n2530,n509,n905);
not gate_2503(n2531,n2530);
and gate_2504(n2532,n2529,n2531);
and gate_2505(n2533,n2515,n2532);
and gate_2506(n2534,n2505,n2533);
not gate_2507(n2535,n2534);
and gate_2508(n2536,n1586,n2535);
not gate_2509(n2537,n2536);
and gate_2510(n2538,n2486,n2537);
and gate_2511(n2539,n2405,n2538);
not gate_2512(n2540,n2539);
and gate_2513(n2541,n32,n2540);
not gate_2514(n2542,n2541);
and gate_2515(n2543,n150,n435);
not gate_2516(n2544,n2543);
and gate_2517(n2545,n1495,n2544);
not gate_2518(n2546,n2545);
and gate_2519(n2547,pi0,n2546);
not gate_2520(n2548,n2547);
and gate_2521(n2549,n1586,n2113);
not gate_2522(n2550,n2549);
and gate_2523(n2551,n2548,n2550);
not gate_2524(n2552,n2551);
and gate_2525(n2553,pi7,n2552);
not gate_2526(n2554,n2553);
and gate_2527(n2555,n30,n1363);
and gate_2528(n2556,n1167,n2555);
not gate_2529(n2557,n2556);
and gate_2530(n2558,n2554,n2557);
not gate_2531(n2559,n2558);
and gate_2532(n2560,n38,n2559);
not gate_2533(n2561,n2560);
and gate_2534(n2562,pi0,n435);
and gate_2535(n2563,n148,n2562);
not gate_2536(n2564,n2563);
and gate_2537(n2565,n2561,n2564);
not gate_2538(n2566,n2565);
and gate_2539(n2567,n33,n2566);
not gate_2540(n2568,n2567);
and gate_2541(n2569,n1543,n1701);
not gate_2542(n2570,n2569);
and gate_2543(n2571,n39,n784);
and gate_2544(n2572,n2570,n2571);
not gate_2545(n2573,n2572);
and gate_2546(n2574,n2568,n2573);
and gate_2547(n2575,n2542,n2574);
and gate_2548(n2576,n2392,n2575);
and gate_2549(n2577,n2156,n2576);
not gate_2550(po06,n2577);
and gate_2551(n2579,n30,pi2);
and gate_2552(n2580,n163,n2579);
not gate_2553(n2581,n2580);
and gate_2554(n2582,pi0,n821);
and gate_2555(n2583,n209,n2582);
not gate_2556(n2584,n2583);
and gate_2557(n2585,n2581,n2584);
not gate_2558(n2586,n2585);
and gate_2559(n2587,n31,n2586);
not gate_2560(n2588,n2587);
and gate_2561(n2589,n821,n2555);
not gate_2562(n2590,n2589);
and gate_2563(n2591,n2588,n2590);
not gate_2564(n2592,n2591);
and gate_2565(n2593,n35,n2592);
not gate_2566(n2594,n2593);
and gate_2567(n2595,n1243,n2100);
not gate_2568(n2596,n2595);
and gate_2569(n2597,n2594,n2596);
not gate_2570(n2598,n2597);
and gate_2571(n2599,n268,n2598);
not gate_2572(n2600,n2599);
and gate_2573(n2601,n819,n2243);
not gate_2574(n2602,n2601);
and gate_2575(n2603,n1730,n2602);
not gate_2576(n2604,n2603);
and gate_2577(n2605,n1282,n2604);
not gate_2578(n2606,n2605);
and gate_2579(n2607,n219,n1586);
not gate_2580(n2608,n2607);
and gate_2581(n2609,pi0,n1202);
and gate_2582(n2610,n224,n2609);
not gate_2583(n2611,n2610);
and gate_2584(n2612,n2608,n2611);
and gate_2585(n2613,n257,n800);
and gate_2586(n2614,pi0,n2613);
not gate_2587(n2615,n2614);
and gate_2588(n2616,n2612,n2615);
not gate_2589(n2617,n2616);
and gate_2590(n2618,pi8,n2617);
not gate_2591(n2619,n2618);
and gate_2592(n2620,n37,n2326);
not gate_2593(n2621,n2620);
and gate_2594(n2622,n69,n257);
not gate_2595(n2623,n2622);
and gate_2596(n2624,n2621,n2623);
not gate_2597(n2625,n2624);
and gate_2598(n2626,pi1,n2625);
not gate_2599(n2627,n2626);
and gate_2600(n2628,n69,n884);
not gate_2601(n2629,n2628);
and gate_2602(n2630,n2627,n2629);
not gate_2603(n2631,n2630);
and gate_2604(n2632,n38,n2631);
not gate_2605(n2633,n2632);
and gate_2606(n2634,n2619,n2633);
not gate_2607(n2635,n2634);
and gate_2608(n2636,n32,n2635);
not gate_2609(n2637,n2636);
and gate_2610(n2638,n1430,n1710);
not gate_2611(n2639,n2638);
and gate_2612(n2640,n388,n1300);
not gate_2613(n2641,n2640);
and gate_2614(n2642,n1975,n2640);
and gate_2615(n2643,n70,n2642);
not gate_2616(n2644,n2643);
and gate_2617(n2645,n2639,n2644);
not gate_2618(n2646,n2645);
and gate_2619(n2647,pi1,n2646);
not gate_2620(n2648,n2647);
and gate_2621(n2649,n30,pi7);
not gate_2622(n2650,n2649);
and gate_2623(n2651,n1842,n2650);
not gate_2624(n2652,n2651);
and gate_2625(n2653,n267,n2652);
and gate_2626(n2654,n192,n2653);
not gate_2627(n2655,n2654);
and gate_2628(n2656,n2648,n2655);
not gate_2629(n2657,n2656);
and gate_2630(n2658,pi2,n2657);
not gate_2631(n2659,n2658);
and gate_2632(n2660,n81,n2243);
not gate_2633(n2661,n2660);
and gate_2634(n2662,n53,n1586);
not gate_2635(n2663,n2662);
and gate_2636(n2664,n2661,n2663);
not gate_2637(n2665,n2664);
and gate_2638(n2666,n142,n2665);
not gate_2639(n2667,n2666);
and gate_2640(n2668,n2659,n2667);
and gate_2641(n2669,n2637,n2668);
and gate_2642(n2670,n2606,n2669);
not gate_2643(n2671,n2670);
and gate_2644(n2672,n35,n2671);
not gate_2645(n2673,n2672);
and gate_2646(n2674,n43,n299);
not gate_2647(n2675,n2674);
and gate_2648(n2676,n1468,n2675);
not gate_2649(n2677,n2676);
and gate_2650(n2678,n30,pi3);
not gate_2651(n2679,n2678);
and gate_2652(n2680,n70,n2679);
not gate_2653(n2681,n2680);
and gate_2654(n2682,n2677,n2681);
not gate_2655(n2683,n2682);
and gate_2656(n2684,pi3,n81);
not gate_2657(n2685,n2684);
and gate_2658(n2686,n33,n53);
not gate_2659(n2687,n2686);
and gate_2660(n2688,n2685,n2687);
not gate_2661(n2689,n2688);
and gate_2662(n2690,n32,n2689);
not gate_2663(n2691,n2690);
and gate_2664(n2692,pi2,n2641);
not gate_2665(n2693,n2692);
and gate_2666(n2694,n2691,n2693);
not gate_2667(n2695,n2694);
and gate_2668(n2696,pi1,n2695);
not gate_2669(n2697,n2696);
and gate_2670(n2698,pi2,pi7);
not gate_2671(n2699,n2698);
and gate_2672(n2700,n749,n2698);
and gate_2673(n2701,n31,n2700);
not gate_2674(n2702,n2701);
and gate_2675(n2703,n2697,n2702);
not gate_2676(n2704,n2703);
and gate_2677(n2705,n30,n2704);
not gate_2678(n2706,n2705);
and gate_2679(n2707,n32,n1489);
not gate_2680(n2708,n2707);
and gate_2681(n2709,n37,n2708);
not gate_2682(n2710,n2709);
and gate_2683(n2711,n32,n39);
not gate_2684(n2712,n2711);
and gate_2685(n2713,n2710,n2712);
not gate_2686(n2714,n2713);
and gate_2687(n2715,n291,n2714);
and gate_2688(n2716,pi0,n2715);
not gate_2689(n2717,n2716);
and gate_2690(n2718,n2706,n2717);
and gate_2691(n2719,n2683,n2718);
not gate_2692(n2720,n2719);
and gate_2693(n2721,pi4,n2720);
not gate_2694(n2722,n2721);
and gate_2695(n2723,pi0,n2689);
not gate_2696(n2724,n2723);
and gate_2697(n2725,n37,n1356);
not gate_2698(n2726,n2725);
and gate_2699(n2727,n40,n2726);
not gate_2700(n2728,n2727);
and gate_2701(n2729,n30,n2728);
not gate_2702(n2730,n2729);
and gate_2703(n2731,n2724,n2730);
not gate_2704(n2732,n2731);
and gate_2705(n2733,n32,n2732);
not gate_2706(n2734,n2733);
and gate_2707(n2735,pi0,n260);
not gate_2708(n2736,n2735);
and gate_2709(n2737,n84,n2736);
not gate_2710(n2738,n2737);
and gate_2711(n2739,n819,n2738);
not gate_2712(n2740,n2739);
and gate_2713(n2741,n2734,n2740);
not gate_2714(n2742,n2741);
and gate_2715(n2743,pi1,n2742);
not gate_2716(n2744,n2743);
and gate_2717(n2745,pi2,n38);
not gate_2718(n2746,n2745);
and gate_2719(n2747,n30,n2745);
not gate_2720(n2748,n2747);
and gate_2721(n2749,n2093,n2641);
not gate_2722(n2750,n2749);
and gate_2723(n2751,n2748,n2750);
not gate_2724(n2752,n2751);
and gate_2725(n2753,n37,n2752);
not gate_2726(n2754,n2753);
and gate_2727(n2755,n1380,n2579);
not gate_2728(n2756,n2755);
and gate_2729(n2757,n2754,n2756);
not gate_2730(n2758,n2757);
and gate_2731(n2759,n31,n2758);
not gate_2732(n2760,n2759);
and gate_2733(n2761,n2744,n2760);
not gate_2734(n2762,n2761);
and gate_2735(n2763,n34,n2762);
not gate_2736(n2764,n2763);
and gate_2737(n2765,n204,n2680);
and gate_2738(n2766,n260,n2765);
and gate_2739(n2767,n1137,n2766);
not gate_2740(n2768,n2767);
and gate_2741(n2769,n2764,n2768);
and gate_2742(n2770,n2722,n2769);
not gate_2743(n2771,n2770);
and gate_2744(n2772,pi5,n2771);
not gate_2745(n2773,n2772);
and gate_2746(n2774,n81,n206);
not gate_2747(n2775,n2774);
and gate_2748(n2776,n636,n1192);
not gate_2749(n2777,n2776);
and gate_2750(n2778,n2775,n2777);
not gate_2751(n2779,n2778);
and gate_2752(n2780,pi1,n2779);
not gate_2753(n2781,n2780);
and gate_2754(n2782,n299,n2686);
not gate_2755(n2783,n2782);
and gate_2756(n2784,n2781,n2783);
not gate_2757(n2785,n2784);
and gate_2758(n2786,pi0,n2785);
not gate_2759(n2787,n2786);
and gate_2760(n2788,n1259,n2774);
not gate_2761(n2789,n2788);
and gate_2762(n2790,n2787,n2789);
and gate_2763(n2791,n2773,n2790);
and gate_2764(n2792,n2673,n2791);
and gate_2765(n2793,n2600,n2792);
not gate_2766(n2794,n2793);
and gate_2767(n2795,pi6,n2794);
not gate_2768(n2796,n2795);
and gate_2769(n2797,n1259,n1754);
not gate_2770(n2798,n2797);
and gate_2771(n2799,n706,n1665);
not gate_2772(n2800,n2799);
and gate_2773(n2801,n2798,n2800);
and gate_2774(n2802,n1542,n1652);
and gate_2775(n2803,pi0,n2802);
not gate_2776(n2804,n2803);
and gate_2777(n2805,n1259,n1634);
not gate_2778(n2806,n2805);
and gate_2779(n2807,n2804,n2806);
and gate_2780(n2808,n1495,n1909);
not gate_2781(n2809,n2808);
and gate_2782(n2810,n30,n2809);
not gate_2783(n2811,n2810);
and gate_2784(n2812,n286,n2243);
not gate_2785(n2813,n2812);
and gate_2786(n2814,n2811,n2813);
not gate_2787(n2815,n2814);
and gate_2788(n2816,pi8,n2815);
not gate_2789(n2817,n2816);
and gate_2790(n2818,n38,n1491);
and gate_2791(n2819,n2395,n2818);
not gate_2792(n2820,n2819);
and gate_2793(n2821,n2817,n2820);
not gate_2794(n2822,n2821);
and gate_2795(n2823,n37,n2822);
not gate_2796(n2824,n2823);
and gate_2797(n2825,n31,pi4);
not gate_2798(n2826,n2825);
and gate_2799(n2827,n455,n2825);
not gate_2800(n2828,n2827);
and gate_2801(n2829,pi1,n99);
not gate_2802(n2830,n2829);
and gate_2803(n2831,n31,n590);
not gate_2804(n2832,n2831);
and gate_2805(n2833,n2830,n2832);
not gate_2806(n2834,n2833);
and gate_2807(n2835,n1762,n2834);
not gate_2808(n2836,n2835);
and gate_2809(n2837,n2828,n2836);
not gate_2810(n2838,n2837);
and gate_2811(n2839,pi7,n2838);
not gate_2812(n2840,n2839);
and gate_2813(n2841,n2824,n2840);
not gate_2814(n2842,n2841);
and gate_2815(n2843,pi2,n2842);
not gate_2816(n2844,n2843);
and gate_2817(n2845,n35,n2735);
not gate_2818(n2846,n2845);
and gate_2819(n2847,n346,n1079);
not gate_2820(n2848,n2847);
and gate_2821(n2849,n2846,n2848);
not gate_2822(n2850,n2849);
and gate_2823(n2851,pi4,n2850);
not gate_2824(n2852,n2851);
and gate_2825(n2853,n38,n44);
not gate_2826(n2854,n2853);
and gate_2827(n2855,n35,n2854);
not gate_2828(n2856,n2855);
and gate_2829(n2857,pi5,n81);
not gate_2830(n2858,n2857);
and gate_2831(n2859,n2856,n2858);
not gate_2832(n2860,n2859);
and gate_2833(n2861,n1552,n2860);
not gate_2834(n2862,n2861);
and gate_2835(n2863,n2852,n2862);
not gate_2836(n2864,n2863);
and gate_2837(n2865,n1145,n2864);
not gate_2838(n2866,n2865);
and gate_2839(n2867,n2844,n2866);
and gate_2840(n2868,n2807,n2867);
and gate_2841(n2869,n2801,n2868);
and gate_2842(n2870,pi2,pi4);
and gate_2843(n2871,n53,n2870);
not gate_2844(n2872,n2871);
and gate_2845(n2873,n889,n1505);
not gate_2846(n2874,n2873);
and gate_2847(n2875,n2872,n2874);
not gate_2848(n2876,n2875);
and gate_2849(n2877,n2396,n2876);
and gate_2850(n2878,n30,n35);
not gate_2851(n2879,n2878);
and gate_2852(n2880,n981,n2879);
and gate_2853(n2881,n2877,n2880);
not gate_2854(n2882,n2881);
and gate_2855(n2883,n2869,n2882);
not gate_2856(n2884,n2883);
and gate_2857(n2885,pi3,n2884);
not gate_2858(n2886,n2885);
and gate_2859(n2887,n888,n1365);
and gate_2860(n2888,n908,n2887);
and gate_2861(n2889,pi0,n2888);
not gate_2862(n2890,n2889);
and gate_2863(n2891,pi1,n37);
not gate_2864(n2892,n2891);
and gate_2865(n2893,pi4,n2892);
not gate_2866(n2894,n2893);
and gate_2867(n2895,n31,n2699);
not gate_2868(n2896,n2895);
and gate_2869(n2897,n2894,n2896);
and gate_2870(n2898,n30,n2897);
not gate_2871(n2899,n2898);
and gate_2872(n2900,n2890,n2899);
not gate_2873(n2901,n2900);
and gate_2874(n2902,pi5,n2901);
not gate_2875(n2903,n2902);
and gate_2876(n2904,pi1,n1975);
and gate_2877(n2905,n30,n2904);
not gate_2878(n2906,n2905);
and gate_2879(n2907,n34,n885);
not gate_2880(n2908,n2907);
and gate_2881(n2909,n2243,n2908);
not gate_2882(n2910,n2909);
and gate_2883(n2911,n2906,n2910);
not gate_2884(n2912,n2911);
and gate_2885(n2913,pi2,n2912);
not gate_2886(n2914,n2913);
and gate_2887(n2915,n907,n970);
and gate_2888(n2916,pi0,n2915);
not gate_2889(n2917,n2916);
and gate_2890(n2918,n2914,n2917);
not gate_2891(n2919,n2918);
and gate_2892(n2920,n35,n2919);
not gate_2893(n2921,n2920);
and gate_2894(n2922,n31,n1324);
and gate_2895(n2923,n2093,n2922);
not gate_2896(n2924,n2923);
and gate_2897(n2925,n2921,n2924);
and gate_2898(n2926,n2903,n2925);
not gate_2899(n2927,n2926);
and gate_2900(n2928,n38,n2927);
not gate_2901(n2929,n2928);
and gate_2902(n2930,n1079,n2895);
not gate_2903(n2931,n2930);
and gate_2904(n2932,n1451,n2931);
not gate_2905(n2933,n2932);
and gate_2906(n2934,pi0,n2933);
not gate_2907(n2935,n2934);
and gate_2908(n2936,pi2,n1179);
not gate_2909(n2937,n2936);
and gate_2910(n2938,n1544,n2937);
not gate_2911(n2939,n2938);
and gate_2912(n2940,n2935,n2939);
not gate_2913(n2941,n2940);
and gate_2914(n2942,pi4,n2941);
not gate_2915(n2943,n2942);
and gate_2916(n2944,n694,n1215);
not gate_2917(n2945,n2944);
and gate_2918(n2946,pi0,pi2);
and gate_2919(n2947,n1078,n2946);
not gate_2920(n2948,n2947);
and gate_2921(n2949,n2945,n2948);
not gate_2922(n2950,n2949);
and gate_2923(n2951,pi1,n2950);
not gate_2924(n2952,n2951);
and gate_2925(n2953,n30,n1577);
not gate_2926(n2954,n2953);
and gate_2927(n2955,n2952,n2954);
not gate_2928(n2956,n2955);
and gate_2929(n2957,n34,n2956);
not gate_2930(n2958,n2957);
and gate_2931(n2959,n2943,n2958);
not gate_2932(n2960,n2959);
and gate_2933(n2961,pi8,n2960);
not gate_2934(n2962,n2961);
and gate_2935(n2963,n1365,n1490);
and gate_2936(n2964,n2244,n2963);
and gate_2937(n2965,n2698,n2964);
not gate_2938(n2966,n2965);
and gate_2939(n2967,n2962,n2966);
and gate_2940(n2968,n2929,n2967);
not gate_2941(n2969,n2968);
and gate_2942(n2970,n33,n2969);
not gate_2943(n2971,n2970);
and gate_2944(n2972,pi0,n1653);
not gate_2945(n2973,n2972);
and gate_2946(n2974,n664,n1506);
and gate_2947(n2975,n2878,n2974);
not gate_2948(n2976,n2975);
and gate_2949(n2977,n2973,n2976);
not gate_2950(n2978,n2977);
and gate_2951(n2979,pi1,n2978);
not gate_2952(n2980,n2979);
and gate_2953(n2981,n813,n1243);
not gate_2954(n2982,n2981);
and gate_2955(n2983,n2980,n2982);
not gate_2956(n2984,n2983);
and gate_2957(n2985,pi7,n2984);
not gate_2958(n2986,n2985);
and gate_2959(n2987,pi0,n299);
and gate_2960(n2988,n43,n509);
and gate_2961(n2989,n2987,n2988);
not gate_2962(n2990,n2989);
and gate_2963(n2991,n2986,n2990);
and gate_2964(n2992,n2971,n2991);
and gate_2965(n2993,n2886,n2992);
not gate_2966(n2994,n2993);
and gate_2967(n2995,n36,n2994);
not gate_2968(n2996,n2995);
and gate_2969(n2997,n30,n953);
and gate_2970(n2998,n53,n608);
and gate_2971(n2999,n2997,n2998);
not gate_2972(n3000,n2999);
and gate_2973(n3001,n897,n1269);
not gate_2974(n3002,n3001);
and gate_2975(n3003,n291,n1273);
not gate_2976(n3004,n3003);
and gate_2977(n3005,n3002,n3004);
not gate_2978(n3006,n3005);
and gate_2979(n3007,n158,n3006);
not gate_2980(n3008,n3007);
and gate_2981(n3009,n3000,n3008);
not gate_2982(n3010,n3009);
and gate_2983(n3011,n32,n3010);
not gate_2984(n3012,n3011);
and gate_2985(n3013,n819,n2395);
and gate_2986(n3014,n43,n277);
and gate_2987(n3015,n3013,n3014);
not gate_2988(n3016,n3015);
and gate_2989(n3017,n3012,n3016);
and gate_2990(n3018,n2996,n3017);
and gate_2991(n3019,n2796,n3018);
not gate_2992(po07,n3019);
and gate_2993(n3021,n299,n560);
not gate_2994(n3022,n3021);
and gate_2995(n3023,n181,n593);
not gate_2996(n3024,n3023);
and gate_2997(n3025,n709,n3024);
not gate_2998(n3026,n3025);
and gate_2999(n3027,n1145,n3026);
not gate_3000(n3028,n3027);
and gate_3001(n3029,n3022,n3028);
not gate_3002(n3030,n3029);
and gate_3003(n3031,n30,n3030);
not gate_3004(n3032,n3031);
and gate_3005(n3033,n1243,n1806);
not gate_3006(n3034,n3033);
and gate_3007(n3035,n3032,n3034);
and gate_3008(n3036,pi8,n229);
not gate_3009(n3037,n3036);
and gate_3010(n3038,n386,n3037);
not gate_3011(n3039,n3038);
and gate_3012(n3040,n180,n3039);
and gate_3013(n3041,pi2,n3040);
not gate_3014(n3042,n3041);
and gate_3015(n3043,pi3,n419);
not gate_3016(n3044,n3043);
and gate_3017(n3045,n1176,n3044);
not gate_3018(n3046,n3045);
and gate_3019(n3047,n3042,n3046);
not gate_3020(n3048,n3047);
and gate_3021(n3049,pi0,n3048);
not gate_3022(n3050,n3049);
and gate_3023(n3051,pi2,n36);
not gate_3024(n3052,n3051);
and gate_3025(n3053,pi3,n1489);
and gate_3026(n3054,n3052,n3053);
not gate_3027(n3055,n3054);
and gate_3028(n3056,n38,n337);
not gate_3029(n3057,n3056);
and gate_3030(n3058,n819,n3057);
not gate_3031(n3059,n3058);
and gate_3032(n3060,n3055,n3059);
not gate_3033(n3061,n3060);
and gate_3034(n3062,n37,n3061);
not gate_3035(n3063,n3062);
and gate_3036(n3064,n104,n1300);
and gate_3037(n3065,n32,n3064);
not gate_3038(n3066,n3065);
and gate_3039(n3067,n3063,n3066);
not gate_3040(n3068,n3067);
and gate_3041(n3069,n30,n3068);
not gate_3042(n3070,n3069);
and gate_3043(n3071,n3050,n3070);
not gate_3044(n3072,n3071);
and gate_3045(n3073,pi5,n3072);
not gate_3046(n3074,n3073);
and gate_3047(n3075,n118,n618);
not gate_3048(n3076,n3075);
and gate_3049(n3077,pi0,n3076);
not gate_3050(n3078,n3077);
and gate_3051(n3079,n43,n135);
not gate_3052(n3080,n3079);
and gate_3053(n3081,n3078,n3080);
not gate_3054(n3082,n3081);
and gate_3055(n3083,n822,n3082);
not gate_3056(n3084,n3083);
and gate_3057(n3085,pi2,pi8);
not gate_3058(n3086,n3085);
and gate_3059(n3087,n32,n748);
not gate_3060(n3088,n3087);
and gate_3061(n3089,n3086,n3088);
not gate_3062(n3090,n3089);
and gate_3063(n3091,n30,n3090);
not gate_3064(n3092,n3091);
and gate_3065(n3093,n387,n2093);
not gate_3066(n3094,n3093);
and gate_3067(n3095,n3092,n3094);
not gate_3068(n3096,n3095);
and gate_3069(n3097,pi7,n3096);
not gate_3070(n3098,n3097);
and gate_3071(n3099,n2582,n2725);
not gate_3072(n3100,n3099);
and gate_3073(n3101,n3098,n3100);
not gate_3074(n3102,n3101);
and gate_3075(n3103,pi6,n3102);
not gate_3076(n3104,n3103);
and gate_3077(n3105,n1380,n2946);
not gate_3078(n3106,n3105);
and gate_3079(n3107,n3104,n3106);
and gate_3080(n3108,n3084,n3107);
not gate_3081(n3109,n3108);
and gate_3082(n3110,n35,n3109);
not gate_3083(n3111,n3110);
and gate_3084(n3112,n3074,n3111);
not gate_3085(n3113,n3112);
and gate_3086(n3114,pi1,n3113);
not gate_3087(n3115,n3114);
and gate_3088(n3116,pi3,n97);
not gate_3089(n3117,n3116);
and gate_3090(n3118,n361,n3117);
and gate_3091(n3119,n33,n1023);
not gate_3092(n3120,n3119);
and gate_3093(n3121,n3118,n3120);
and gate_3094(n3122,n35,n3121);
not gate_3095(n3123,n3122);
and gate_3096(n3124,n46,n659);
not gate_3097(n3125,n3124);
and gate_3098(n3126,pi3,n3125);
not gate_3099(n3127,n3126);
and gate_3100(n3128,n66,n3127);
not gate_3101(n3129,n3128);
and gate_3102(n3130,pi5,n3129);
not gate_3103(n3131,n3130);
and gate_3104(n3132,n3123,n3131);
not gate_3105(n3133,n3132);
and gate_3106(n3134,pi0,n3133);
not gate_3107(n3135,n3134);
and gate_3108(n3136,n35,n883);
not gate_3109(n3137,n3136);
and gate_3110(n3138,n37,n82);
not gate_3111(n3139,n3138);
and gate_3112(n3140,n150,n3139);
not gate_3113(n3141,n3140);
and gate_3114(n3142,n3137,n3141);
not gate_3115(n3143,n3142);
and gate_3116(n3144,n1692,n3143);
not gate_3117(n3145,n3144);
and gate_3118(n3146,n3135,n3145);
not gate_3119(n3147,n3146);
and gate_3120(n3148,pi2,n3147);
not gate_3121(n3149,n3148);
and gate_3122(n3150,n337,n906);
not gate_3123(n3151,n3150);
and gate_3124(n3152,n33,n3151);
not gate_3125(n3153,n3152);
and gate_3126(n3154,n39,n309);
not gate_3127(n3155,n3154);
and gate_3128(n3156,n3153,n3155);
not gate_3129(n3157,n3156);
and gate_3130(n3158,n35,n3157);
not gate_3131(n3159,n3158);
and gate_3132(n3160,n337,n585);
not gate_3133(n3161,n3160);
and gate_3134(n3162,n114,n3161);
not gate_3135(n3163,n3162);
and gate_3136(n3164,n3159,n3163);
not gate_3137(n3165,n3164);
and gate_3138(n3166,n32,n3165);
not gate_3139(n3167,n3166);
and gate_3140(n3168,n177,n593);
and gate_3141(n3169,n219,n3168);
not gate_3142(n3170,n3169);
and gate_3143(n3171,n3167,n3170);
not gate_3144(n3172,n3171);
and gate_3145(n3173,pi0,n3172);
not gate_3146(n3174,n3173);
and gate_3147(n3175,n3149,n3174);
not gate_3148(n3176,n3175);
and gate_3149(n3177,n31,n3176);
not gate_3150(n3178,n3177);
and gate_3151(n3179,pi8,n1006);
and gate_3152(n3180,n224,n3179);
and gate_3153(n3181,pi0,n3180);
not gate_3154(n3182,n3181);
and gate_3155(n3183,n131,n1692);
not gate_3156(n3184,n3183);
and gate_3157(n3185,n3182,n3184);
not gate_3158(n3186,n3185);
and gate_3159(n3187,n36,n3186);
not gate_3160(n3188,n3187);
and gate_3161(n3189,n30,n239);
and gate_3162(n3190,n117,n3189);
not gate_3163(n3191,n3190);
and gate_3164(n3192,n3188,n3191);
not gate_3165(n3193,n3192);
and gate_3166(n3194,pi2,n3193);
not gate_3167(n3195,n3194);
and gate_3168(n3196,pi0,n1154);
and gate_3169(n3197,n43,n146);
and gate_3170(n3198,n3196,n3197);
not gate_3171(n3199,n3198);
and gate_3172(n3200,n3195,n3199);
and gate_3173(n3201,n3178,n3200);
and gate_3174(n3202,n3115,n3201);
and gate_3175(n3203,n3035,n3202);
not gate_3176(n3204,n3203);
and gate_3177(n3205,n34,n3204);
not gate_3178(n3206,n3205);
and gate_3179(n3207,n118,n1822);
not gate_3180(n3208,n3207);
and gate_3181(n3209,n33,n3208);
not gate_3182(n3210,n3209);
and gate_3183(n3211,n53,n175);
not gate_3184(n3212,n3211);
and gate_3185(n3213,n66,n333);
not gate_3186(n3214,n3213);
and gate_3187(n3215,n239,n3214);
not gate_3188(n3216,n3215);
and gate_3189(n3217,n3212,n3216);
and gate_3190(n3218,n3210,n3217);
not gate_3191(n3219,n3218);
and gate_3192(n3220,pi2,n3219);
not gate_3193(n3221,n3220);
and gate_3194(n3222,pi5,n52);
not gate_3195(n3223,n3222);
and gate_3196(n3224,pi7,n310);
and gate_3197(n3225,n3223,n3224);
not gate_3198(n3226,n3225);
and gate_3199(n3227,n1955,n3226);
not gate_3200(n3228,n3227);
and gate_3201(n3229,pi8,n3228);
not gate_3202(n3230,n3229);
and gate_3203(n3231,pi5,n228);
not gate_3204(n3232,n3231);
and gate_3205(n3233,n37,n226);
not gate_3206(n3234,n3233);
and gate_3207(n3235,n3232,n3234);
and gate_3208(n3236,n38,n3235);
not gate_3209(n3237,n3236);
and gate_3210(n3238,n242,n3237);
and gate_3211(n3239,n3230,n3238);
not gate_3212(n3240,n3239);
and gate_3213(n3241,n32,n3240);
not gate_3214(n3242,n3241);
and gate_3215(n3243,n3221,n3242);
not gate_3216(n3244,n3243);
and gate_3217(n3245,pi0,n3244);
not gate_3218(n3246,n3245);
and gate_3219(n3247,n590,n1154);
not gate_3220(n3248,n3247);
and gate_3221(n3249,n32,n99);
not gate_3222(n3250,n3249);
and gate_3223(n3251,n1578,n3250);
not gate_3224(n3252,n3251);
and gate_3225(n3253,pi3,n3251);
not gate_3226(n3254,n3253);
and gate_3227(n3255,n3248,n3254);
not gate_3228(n3256,n3255);
and gate_3229(n3257,pi7,n3256);
not gate_3230(n3258,n3257);
and gate_3231(n3259,pi3,n3252);
not gate_3232(n3260,n3259);
and gate_3233(n3261,n819,n2292);
not gate_3234(n3262,n3261);
and gate_3235(n3263,n3260,n3262);
not gate_3236(n3264,n3263);
and gate_3237(n3265,n37,n3264);
not gate_3238(n3266,n3265);
and gate_3239(n3267,n3258,n3266);
not gate_3240(n3268,n3267);
and gate_3241(n3269,n30,n3268);
not gate_3242(n3270,n3269);
and gate_3243(n3271,n81,n217);
not gate_3244(n3272,n3271);
and gate_3245(n3273,n3270,n3272);
not gate_3246(n3274,n3273);
and gate_3247(n3275,pi6,n3274);
not gate_3248(n3276,n3275);
and gate_3249(n3277,n32,n711);
not gate_3250(n3278,n3277);
and gate_3251(n3279,n561,n3278);
not gate_3252(n3280,n3279);
and gate_3253(n3281,n30,n3280);
not gate_3254(n3282,n3281);
and gate_3255(n3283,n39,n1063);
not gate_3256(n3284,n3283);
and gate_3257(n3285,n3282,n3284);
not gate_3258(n3286,n3285);
and gate_3259(n3287,n33,n3286);
not gate_3260(n3288,n3287);
and gate_3261(n3289,pi2,n1128);
not gate_3262(n3290,n3289);
and gate_3263(n3291,pi2,n3290);
not gate_3264(n3292,n3291);
and gate_3265(n3293,n1299,n3292);
and gate_3266(n3294,n30,n3293);
not gate_3267(n3295,n3294);
and gate_3268(n3296,n3288,n3295);
not gate_3269(n3297,n3296);
and gate_3270(n3298,n36,n3297);
not gate_3271(n3299,n3298);
and gate_3272(n3300,n3276,n3299);
and gate_3273(n3301,n3246,n3300);
not gate_3274(n3302,n3301);
and gate_3275(n3303,pi1,n3302);
not gate_3276(n3304,n3303);
and gate_3277(n3305,pi0,n421);
not gate_3278(n3306,n3305);
and gate_3279(n3307,n30,n418);
not gate_3280(n3308,n3307);
and gate_3281(n3309,n3306,n3308);
not gate_3282(n3310,n3309);
and gate_3283(n3311,pi5,n3310);
not gate_3284(n3312,n3311);
and gate_3285(n3313,n30,n99);
not gate_3286(n3314,n3313);
and gate_3287(n3315,n3312,n3314);
not gate_3288(n3316,n3315);
and gate_3289(n3317,pi3,n3316);
not gate_3290(n3318,n3317);
and gate_3291(n3319,n147,n151);
not gate_3292(n3320,n3319);
and gate_3293(n3321,n2147,n3319);
not gate_3294(n3322,n3321);
and gate_3295(n3323,n748,n3322);
not gate_3296(n3324,n3323);
and gate_3297(n3325,n3318,n3324);
not gate_3298(n3326,n3325);
and gate_3299(n3327,pi2,n3326);
not gate_3300(n3328,n3327);
and gate_3301(n3329,n51,n592);
not gate_3302(n3330,n3329);
and gate_3303(n3331,n52,n593);
not gate_3304(n3332,n3331);
and gate_3305(n3333,n3330,n3332);
not gate_3306(n3334,n3333);
and gate_3307(n3335,n520,n3334);
and gate_3308(n3336,n32,n3335);
not gate_3309(n3337,n3336);
and gate_3310(n3338,n217,n418);
not gate_3311(n3339,n3338);
and gate_3312(n3340,n3337,n3339);
not gate_3313(n3341,n3340);
and gate_3314(n3342,pi0,n3341);
not gate_3315(n3343,n3342);
and gate_3316(n3344,n3328,n3343);
not gate_3317(n3345,n3344);
and gate_3318(n3346,n37,n3345);
not gate_3319(n3347,n3346);
and gate_3320(n3348,pi0,n226);
not gate_3321(n3349,n3348);
and gate_3322(n3350,n88,n228);
and gate_3323(n3351,n3349,n3350);
and gate_3324(n3352,n38,n3351);
not gate_3325(n3353,n3352);
and gate_3326(n3354,n35,n2198);
not gate_3327(n3355,n3354);
and gate_3328(n3356,n3308,n3355);
not gate_3329(n3357,n3356);
and gate_3330(n3358,n2879,n3357);
not gate_3331(n3359,n3358);
and gate_3332(n3360,n3353,n3359);
not gate_3333(n3361,n3360);
and gate_3334(n3362,pi2,n3361);
not gate_3335(n3363,n3362);
and gate_3336(n3364,n35,n421);
not gate_3337(n3365,n3364);
and gate_3338(n3366,n1872,n3365);
not gate_3339(n3367,n3366);
and gate_3340(n3368,n33,n3367);
not gate_3341(n3369,n3368);
and gate_3342(n3370,n52,n455);
not gate_3343(n3371,n3370);
and gate_3344(n3372,n3369,n3371);
not gate_3345(n3373,n3372);
and gate_3346(n3374,n2093,n3373);
not gate_3347(n3375,n3374);
and gate_3348(n3376,n3363,n3375);
not gate_3349(n3377,n3376);
and gate_3350(n3378,pi7,n3377);
not gate_3351(n3379,n3378);
and gate_3352(n3380,n30,n819);
and gate_3353(n3381,n528,n3380);
not gate_3354(n3382,n3381);
and gate_3355(n3383,n3379,n3382);
and gate_3356(n3384,n3347,n3383);
not gate_3357(n3385,n3384);
and gate_3358(n3386,n31,n3385);
not gate_3359(n3387,n3386);
and gate_3360(n3388,n3304,n3387);
not gate_3361(n3389,n3388);
and gate_3362(n3390,pi4,n3389);
not gate_3363(n3391,n3390);
and gate_3364(n3392,n560,n1710);
not gate_3365(n3393,n3392);
and gate_3366(n3394,n130,n695);
not gate_3367(n3395,n3394);
and gate_3368(n3396,n1692,n3395);
not gate_3369(n3397,n3396);
and gate_3370(n3398,n3393,n3397);
not gate_3371(n3399,n3398);
and gate_3372(n3400,n32,n3399);
not gate_3373(n3401,n3400);
and gate_3374(n3402,n957,n3380);
not gate_3375(n3403,n3402);
and gate_3376(n3404,n3401,n3403);
not gate_3377(n3405,n3404);
and gate_3378(n3406,n1048,n3405);
not gate_3379(n3407,n3406);
and gate_3380(n3408,n3391,n3407);
and gate_3381(n3409,n3206,n3408);
not gate_3382(po08,n3409);
and gate_3383(n3411,n1259,n2988);
not gate_3384(n3412,n3411);
and gate_3385(n3413,n81,n2870);
not gate_3386(n3414,n3413);
and gate_3387(n3415,n53,n907);
not gate_3388(n3416,n3415);
and gate_3389(n3417,n3414,n3416);
not gate_3390(n3418,n3417);
and gate_3391(n3419,pi0,n3418);
not gate_3392(n3420,n3419);
and gate_3393(n3421,n34,n43);
not gate_3394(n3422,n3421);
and gate_3395(n3423,n1327,n3422);
not gate_3396(n3424,n3423);
and gate_3397(n3425,n2579,n3424);
not gate_3398(n3426,n3425);
and gate_3399(n3427,n3420,n3426);
not gate_3400(n3428,n3427);
and gate_3401(n3429,n1542,n3428);
not gate_3402(n3430,n3429);
and gate_3403(n3431,n3412,n3430);
not gate_3404(n3432,n3431);
and gate_3405(n3433,n230,n3432);
not gate_3406(n3434,n3433);
and gate_3407(n3435,n32,pi6);
not gate_3408(n3436,n3435);
and gate_3409(n3437,n3052,n3436);
not gate_3410(n3438,n3437);
and gate_3411(n3439,n1365,n2134);
and gate_3412(n3440,n3438,n3439);
not gate_3413(n3441,n3440);
and gate_3414(n3442,n30,n3441);
not gate_3415(n3443,n3442);
and gate_3416(n3444,n2651,n3443);
and gate_3417(n3445,n627,n785);
not gate_3418(n3446,n3445);
and gate_3419(n3447,n1186,n1251);
and gate_3420(n3448,n3446,n3447);
not gate_3421(n3449,n3448);
and gate_3422(n3450,pi0,n3449);
not gate_3423(n3451,n3450);
and gate_3424(n3452,n3444,n3451);
and gate_3425(n3453,pi3,n3452);
not gate_3426(n3454,n3453);
and gate_3427(n3455,n30,n3435);
not gate_3428(n3456,n3455);
and gate_3429(n3457,n191,n2946);
not gate_3430(n3458,n3457);
and gate_3431(n3459,n3456,n3458);
not gate_3432(n3460,n3459);
and gate_3433(n3461,n34,n3460);
not gate_3434(n3462,n3461);
and gate_3435(n3463,n626,n2937);
and gate_3436(n3464,n30,n3463);
not gate_3437(n3465,n3464);
and gate_3438(n3466,n3462,n3465);
not gate_3439(n3467,n3466);
and gate_3440(n3468,n897,n3467);
not gate_3441(n3469,n3468);
and gate_3442(n3470,n3454,n3469);
and gate_3443(n3471,pi0,n1505);
not gate_3444(n3472,n3471);
and gate_3445(n3473,n2748,n3472);
not gate_3446(n3474,n3473);
and gate_3447(n3475,n205,n3474);
not gate_3448(n3476,n3475);
and gate_3449(n3477,n30,n820);
not gate_3450(n3478,n3477);
and gate_3451(n3479,n205,n1193);
not gate_3452(n3480,n3479);
and gate_3453(n3481,n3478,n3480);
and gate_3454(n3482,pi8,n3481);
not gate_3455(n3483,n3482);
and gate_3456(n3484,n3476,n3483);
not gate_3457(n3485,n3484);
and gate_3458(n3486,pi6,n3485);
not gate_3459(n3487,n3486);
and gate_3460(n3488,n38,n1476);
not gate_3461(n3489,n3488);
and gate_3462(n3490,pi3,n3489);
not gate_3463(n3491,n3490);
and gate_3464(n3492,n32,n1177);
not gate_3465(n3493,n3492);
and gate_3466(n3494,n748,n3493);
not gate_3467(n3495,n3494);
and gate_3468(n3496,n3491,n3495);
not gate_3469(n3497,n3496);
and gate_3470(n3498,n137,n3497);
not gate_3471(n3499,n3498);
and gate_3472(n3500,n3487,n3499);
not gate_3473(n3501,n3500);
and gate_3474(n3502,n31,n3501);
not gate_3475(n3503,n3502);
and gate_3476(n3504,n30,n419);
not gate_3477(n3505,n3504);
and gate_3478(n3506,n1489,n3086);
not gate_3479(n3507,n3506);
and gate_3480(n3508,n337,n3507);
not gate_3481(n3509,n3508);
and gate_3482(n3510,n3505,n3509);
and gate_3483(n3511,n37,n3510);
not gate_3484(n3512,n3511);
and gate_3485(n3513,n135,n2746);
not gate_3486(n3514,n3513);
and gate_3487(n3515,n1919,n3514);
not gate_3488(n3516,n3515);
and gate_3489(n3517,pi7,n3516);
not gate_3490(n3518,n3517);
and gate_3491(n3519,n3512,n3518);
not gate_3492(n3520,n3519);
and gate_3493(n3521,pi3,n3520);
not gate_3494(n3522,n3521);
and gate_3495(n3523,n40,n182);
not gate_3496(n3524,n3523);
and gate_3497(n3525,pi0,n3524);
not gate_3498(n3526,n3525);
and gate_3499(n3527,n3308,n3526);
not gate_3500(n3528,n3527);
and gate_3501(n3529,n32,n3528);
not gate_3502(n3530,n3529);
and gate_3503(n3531,pi6,n2652);
not gate_3504(n3532,n3531);
and gate_3505(n3533,n180,n3532);
not gate_3506(n3534,n3533);
and gate_3507(n3535,n3085,n3534);
not gate_3508(n3536,n3535);
and gate_3509(n3537,n3530,n3536);
not gate_3510(n3538,n3537);
and gate_3511(n3539,n33,n3538);
not gate_3512(n3540,n3539);
and gate_3513(n3541,n41,n2579);
not gate_3514(n3542,n3541);
and gate_3515(n3543,n3540,n3542);
and gate_3516(n3544,n3522,n3543);
not gate_3517(n3545,n3544);
and gate_3518(n3546,pi1,n3545);
not gate_3519(n3547,n3546);
and gate_3520(n3548,n3503,n3547);
not gate_3521(n3549,n3548);
and gate_3522(n3550,pi4,n3549);
not gate_3523(n3551,n3550);
and gate_3524(n3552,pi8,n1049);
not gate_3525(n3553,n3552);
and gate_3526(n3554,n97,n3553);
not gate_3527(n3555,n3554);
and gate_3528(n3556,n98,n3552);
not gate_3529(n3557,n3556);
and gate_3530(n3558,n3555,n3557);
and gate_3531(n3559,pi0,n3558);
not gate_3532(n3560,n3559);
and gate_3533(n3561,n31,n333);
not gate_3534(n3562,n3561);
and gate_3535(n3563,n37,n337);
not gate_3536(n3564,n3563);
and gate_3537(n3565,n3562,n3564);
and gate_3538(n3566,n30,n3565);
not gate_3539(n3567,n3566);
and gate_3540(n3568,n3560,n3567);
not gate_3541(n3569,n3568);
and gate_3542(n3570,pi3,n3569);
not gate_3543(n3571,n3570);
and gate_3544(n3572,pi1,n1528);
not gate_3545(n3573,n3572);
and gate_3546(n3574,pi0,n3573);
not gate_3547(n3575,n3574);
and gate_3548(n3576,n1537,n3575);
not gate_3549(n3577,n3576);
and gate_3550(n3578,n37,n3577);
not gate_3551(n3579,n3578);
and gate_3552(n3580,n314,n3579);
not gate_3553(n3581,n3580);
and gate_3554(n3582,pi6,n3581);
not gate_3555(n3583,n3582);
and gate_3556(n3584,n314,n337);
not gate_3557(n3585,n3584);
and gate_3558(n3586,n250,n3585);
and gate_3559(n3587,pi7,n3586);
not gate_3560(n3588,n3587);
and gate_3561(n3589,n3583,n3588);
not gate_3562(n3590,n3589);
and gate_3563(n3591,n33,n3590);
not gate_3564(n3592,n3591);
and gate_3565(n3593,n3571,n3592);
not gate_3566(n3594,n3593);
and gate_3567(n3595,pi2,n3594);
not gate_3568(n3596,n3595);
and gate_3569(n3597,n30,n37);
not gate_3570(n3598,n3597);
and gate_3571(n3599,n38,n3598);
not gate_3572(n3600,n3599);
and gate_3573(n3601,n140,n1842);
not gate_3574(n3602,n3601);
and gate_3575(n3603,n3600,n3602);
and gate_3576(n3604,pi1,n3603);
not gate_3577(n3605,n3604);
and gate_3578(n3606,n2236,n3605);
not gate_3579(n3607,n3606);
and gate_3580(n3608,pi3,n3607);
not gate_3581(n3609,n3608);
and gate_3582(n3610,n31,n3151);
not gate_3583(n3611,n3610);
and gate_3584(n3612,n190,n2892);
not gate_3585(n3613,n3612);
and gate_3586(n3614,n38,n3613);
not gate_3587(n3615,n3614);
and gate_3588(n3616,n3611,n3615);
not gate_3589(n3617,n3616);
and gate_3590(n3618,n69,n3617);
not gate_3591(n3619,n3618);
and gate_3592(n3620,n3609,n3619);
not gate_3593(n3621,n3620);
and gate_3594(n3622,n32,n3621);
not gate_3595(n3623,n3622);
and gate_3596(n3624,n584,n801);
not gate_3597(n3625,n3624);
and gate_3598(n3626,n3623,n3625);
and gate_3599(n3627,n3596,n3626);
not gate_3600(n3628,n3627);
and gate_3601(n3629,n34,n3628);
not gate_3602(n3630,n3629);
and gate_3603(n3631,n84,n2687);
not gate_3604(n3632,n3631);
and gate_3605(n3633,pi6,n3632);
and gate_3606(n3634,n299,n3633);
not gate_3607(n3635,n3634);
and gate_3608(n3636,n3630,n3635);
and gate_3609(n3637,n3551,n3636);
and gate_3610(n3638,n3470,n3637);
not gate_3611(n3639,n3638);
and gate_3612(n3640,n35,n3639);
not gate_3613(n3641,n3640);
and gate_3614(n3642,n786,n2395);
not gate_3615(n3643,n3642);
and gate_3616(n3644,pi1,n424);
not gate_3617(n3645,n3644);
and gate_3618(n3646,n2210,n3645);
not gate_3619(n3647,n3646);
and gate_3620(n3648,n2678,n3647);
not gate_3621(n3649,n3648);
and gate_3622(n3650,n3643,n3649);
and gate_3623(n3651,n30,n3446);
not gate_3624(n3652,n3651);
and gate_3625(n3653,n2337,n3652);
not gate_3626(n3654,n3653);
and gate_3627(n3655,pi1,n3654);
not gate_3628(n3656,n3655);
and gate_3629(n3657,pi6,n359);
not gate_3630(n3658,n3657);
and gate_3631(n3659,pi4,n3658);
not gate_3632(n3660,n3659);
and gate_3633(n3661,n1265,n3660);
not gate_3634(n3662,n3661);
and gate_3635(n3663,n2243,n3662);
not gate_3636(n3664,n3663);
and gate_3637(n3665,n3656,n3664);
not gate_3638(n3666,n3665);
and gate_3639(n3667,pi3,n3666);
not gate_3640(n3668,n3667);
and gate_3641(n3669,pi0,n336);
not gate_3642(n3670,n3669);
and gate_3643(n3671,pi4,n333);
not gate_3644(n3672,n3671);
and gate_3645(n3673,n3670,n3672);
not gate_3646(n3674,n3673);
and gate_3647(n3675,n31,n3674);
not gate_3648(n3676,n3675);
and gate_3649(n3677,pi4,n418);
not gate_3650(n3678,n3677);
and gate_3651(n3679,n1586,n3677);
not gate_3652(n3680,n3679);
and gate_3653(n3681,n3676,n3680);
not gate_3654(n3682,n3681);
and gate_3655(n3683,n33,n3682);
not gate_3656(n3684,n3683);
and gate_3657(n3685,n3668,n3684);
and gate_3658(n3686,n3650,n3685);
not gate_3659(n3687,n3686);
and gate_3660(n3688,n37,n3687);
not gate_3661(n3689,n3688);
and gate_3662(n3690,n373,n1537);
and gate_3663(n3691,n480,n2398);
not gate_3664(n3692,n3691);
and gate_3665(n3693,n3690,n3692);
not gate_3666(n3694,n3693);
and gate_3667(n3695,pi3,n3694);
not gate_3668(n3696,n3695);
and gate_3669(n3697,n314,n1366);
not gate_3670(n3698,n3697);
and gate_3671(n3699,n966,n3698);
and gate_3672(n3700,n33,n3699);
not gate_3673(n3701,n3700);
and gate_3674(n3702,n3696,n3701);
not gate_3675(n3703,n3702);
and gate_3676(n3704,n36,n3703);
not gate_3677(n3705,n3704);
and gate_3678(n3706,n33,n662);
and gate_3679(n3707,n2395,n3706);
not gate_3680(n3708,n3707);
and gate_3681(n3709,n208,n436);
and gate_3682(n3710,n346,n3709);
not gate_3683(n3711,n3710);
and gate_3684(n3712,n3708,n3711);
not gate_3685(n3713,n3712);
and gate_3686(n3714,pi6,n3713);
not gate_3687(n3715,n3714);
and gate_3688(n3716,n3705,n3715);
not gate_3689(n3717,n3716);
and gate_3690(n3718,pi7,n3717);
not gate_3691(n3719,n3718);
and gate_3692(n3720,n30,n897);
and gate_3693(n3721,n412,n3720);
not gate_3694(n3722,n3721);
and gate_3695(n3723,n3719,n3722);
and gate_3696(n3724,n3689,n3723);
not gate_3697(n3725,n3724);
and gate_3698(n3726,pi5,n3725);
not gate_3699(n3727,n3726);
and gate_3700(n3728,n358,n869);
not gate_3701(n3729,n3728);
and gate_3702(n3730,n1158,n3729);
not gate_3703(n3731,n3730);
and gate_3704(n3732,pi0,n3731);
not gate_3705(n3733,n3732);
and gate_3706(n3734,n30,n869);
and gate_3707(n3735,n905,n3734);
not gate_3708(n3736,n3735);
and gate_3709(n3737,n3733,n3736);
not gate_3710(n3738,n3737);
and gate_3711(n3739,pi3,n3738);
not gate_3712(n3740,n3739);
and gate_3713(n3741,n30,n799);
and gate_3714(n3742,n628,n3741);
not gate_3715(n3743,n3742);
and gate_3716(n3744,n3740,n3743);
and gate_3717(n3745,n3727,n3744);
not gate_3718(n3746,n3745);
and gate_3719(n3747,pi2,n3746);
not gate_3720(n3748,n3747);
and gate_3721(n3749,n34,n203);
and gate_3722(n3750,n105,n3749);
not gate_3723(n3751,n3750);
and gate_3724(n3752,n2123,n3751);
not gate_3725(n3753,n3752);
and gate_3726(n3754,n31,n3753);
not gate_3727(n3755,n3754);
and gate_3728(n3756,n186,n645);
not gate_3729(n3757,n3756);
and gate_3730(n3758,n953,n3757);
not gate_3731(n3759,n3758);
and gate_3732(n3760,n3755,n3759);
not gate_3733(n3761,n3760);
and gate_3734(n3762,n38,n3761);
not gate_3735(n3763,n3762);
and gate_3736(n3764,n1702,n3445);
and gate_3737(n3765,n1975,n3764);
and gate_3738(n3766,n31,n3765);
not gate_3739(n3767,n3766);
and gate_3740(n3768,n309,n2894);
not gate_3741(n3769,n3768);
and gate_3742(n3770,n3767,n3769);
not gate_3743(n3771,n3770);
and gate_3744(n3772,pi8,n3771);
not gate_3745(n3773,n3772);
and gate_3746(n3774,n3763,n3773);
not gate_3747(n3775,n3774);
and gate_3748(n3776,pi0,n3775);
not gate_3749(n3777,n3776);
and gate_3750(n3778,pi4,n312);
not gate_3751(n3779,n3778);
and gate_3752(n3780,n143,n3779);
not gate_3753(n3781,n3780);
and gate_3754(n3782,n260,n3781);
not gate_3755(n3783,n3782);
and gate_3756(n3784,pi3,n784);
not gate_3757(n3785,n3784);
and gate_3758(n3786,n224,n626);
not gate_3759(n3787,n3786);
and gate_3760(n3788,n3785,n3787);
not gate_3761(n3789,n3788);
and gate_3762(n3790,n38,n3789);
not gate_3763(n3791,n3790);
and gate_3764(n3792,pi3,n1269);
not gate_3765(n3793,n3792);
and gate_3766(n3794,n3791,n3793);
and gate_3767(n3795,n3783,n3794);
not gate_3768(n3796,n3795);
and gate_3769(n3797,n1586,n3796);
not gate_3770(n3798,n3797);
and gate_3771(n3799,n3777,n3798);
not gate_3772(n3800,n3799);
and gate_3773(n3801,pi5,n3800);
not gate_3774(n3802,n3801);
and gate_3775(n3803,pi1,n626);
not gate_3776(n3804,n3803);
and gate_3777(n3805,n179,n435);
not gate_3778(n3806,n3805);
and gate_3779(n3807,n3804,n3806);
not gate_3780(n3808,n3807);
and gate_3781(n3809,n387,n3808);
and gate_3782(n3810,pi0,n3809);
not gate_3783(n3811,n3810);
and gate_3784(n3812,n3802,n3811);
not gate_3785(n3813,n3812);
and gate_3786(n3814,n32,n3813);
not gate_3787(n3815,n3814);
and gate_3788(n3816,n104,n2562);
not gate_3789(n3817,n3816);
and gate_3790(n3818,n97,n2555);
not gate_3791(n3819,n3818);
and gate_3792(n3820,n3817,n3819);
not gate_3793(n3821,n3820);
and gate_3794(n3822,n33,n590);
and gate_3795(n3823,n3821,n3822);
not gate_3796(n3824,n3823);
and gate_3797(n3825,n3815,n3824);
and gate_3798(n3826,n3748,n3825);
and gate_3799(n3827,n3641,n3826);
and gate_3800(n3828,n3434,n3827);
not gate_3801(po09,n3828);
and gate_3802(n3830,n30,n582);
not gate_3803(n3831,n3830);
and gate_3804(n3832,n278,n1587);
not gate_3805(n3833,n3832);
and gate_3806(n3834,n3831,n3833);
and gate_3807(n3835,n33,n3834);
not gate_3808(n3836,n3835);
and gate_3809(n3837,pi3,n608);
and gate_3810(n3838,n2243,n3837);
not gate_3811(n3839,n3838);
and gate_3812(n3840,n3836,n3839);
not gate_3813(n3841,n3840);
and gate_3814(n3842,n32,n3841);
not gate_3815(n3843,n3842);
and gate_3816(n3844,n33,n285);
and gate_3817(n3845,n1259,n3844);
not gate_3818(n3846,n3845);
and gate_3819(n3847,n3843,n3846);
not gate_3820(n3848,n3847);
and gate_3821(n3849,n260,n3848);
not gate_3822(n3850,n3849);
and gate_3823(n3851,n34,n706);
not gate_3824(n3852,n3851);
and gate_3825(n3853,n1755,n3852);
not gate_3826(n3854,n3853);
and gate_3827(n3855,n1586,n2745);
not gate_3828(n3856,n3855);
and gate_3829(n3857,n344,n1243);
not gate_3830(n3858,n3857);
and gate_3831(n3859,n3856,n3858);
not gate_3832(n3860,n3859);
and gate_3833(n3861,n3854,n3860);
not gate_3834(n3862,n3861);
and gate_3835(n3863,pi8,n821);
not gate_3836(n3864,n3863);
and gate_3837(n3865,n38,n822);
not gate_3838(n3866,n3865);
and gate_3839(n3867,n3864,n3866);
not gate_3840(n3868,n3867);
and gate_3841(n3869,n1254,n3868);
and gate_3842(n3870,pi7,n3869);
not gate_3843(n3871,n3870);
and gate_3844(n3872,n82,n591);
not gate_3845(n3873,n3872);
and gate_3846(n3874,n218,n3873);
and gate_3847(n3875,pi2,n3874);
not gate_3848(n3876,n3875);
and gate_3849(n3877,n3871,n3876);
not gate_3850(n3878,n3877);
and gate_3851(n3879,n34,n3878);
not gate_3852(n3880,n3879);
and gate_3853(n3881,n1180,n1489);
and gate_3854(n3882,n1193,n3881);
and gate_3855(n3883,pi5,n3882);
not gate_3856(n3884,n3883);
and gate_3857(n3885,pi2,n387);
and gate_3858(n3886,n707,n3885);
not gate_3859(n3887,n3886);
and gate_3860(n3888,n3884,n3887);
and gate_3861(n3889,n821,n2640);
and gate_3862(n3890,n1181,n3889);
not gate_3863(n3891,n3890);
and gate_3864(n3892,n3888,n3891);
not gate_3865(n3893,n3892);
and gate_3866(n3894,pi4,n3893);
not gate_3867(n3895,n3894);
and gate_3868(n3896,n3880,n3895);
not gate_3869(n3897,n3896);
and gate_3870(n3898,pi0,n3897);
not gate_3871(n3899,n3898);
and gate_3872(n3900,n563,n1327);
not gate_3873(n3901,n3900);
and gate_3874(n3902,n35,n3901);
not gate_3875(n3903,n3902);
and gate_3876(n3904,n53,n509);
not gate_3877(n3905,n3904);
and gate_3878(n3906,n3903,n3905);
not gate_3879(n3907,n3906);
and gate_3880(n3908,n33,n3907);
not gate_3881(n3909,n3908);
and gate_3882(n3910,n34,n3395);
not gate_3883(n3911,n3910);
and gate_3884(n3912,n81,n277);
not gate_3885(n3913,n3912);
and gate_3886(n3914,n3911,n3913);
not gate_3887(n3915,n3914);
and gate_3888(n3916,pi3,n3915);
not gate_3889(n3917,n3916);
and gate_3890(n3918,n3909,n3917);
not gate_3891(n3919,n3918);
and gate_3892(n3920,n32,n3919);
not gate_3893(n3921,n3920);
and gate_3894(n3922,n209,n3085);
not gate_3895(n3923,n3922);
and gate_3896(n3924,n929,n3923);
not gate_3897(n3925,n3924);
and gate_3898(n3926,n37,n3925);
not gate_3899(n3927,n3926);
and gate_3900(n3928,n53,n142);
not gate_3901(n3929,n3928);
and gate_3902(n3930,n3927,n3929);
not gate_3903(n3931,n3930);
and gate_3904(n3932,n35,n3931);
not gate_3905(n3933,n3932);
and gate_3906(n3934,n78,n163);
not gate_3907(n3935,n3934);
and gate_3908(n3936,n1937,n3935);
not gate_3909(n3937,n3936);
and gate_3910(n3938,n1577,n3937);
not gate_3911(n3939,n3938);
and gate_3912(n3940,n3933,n3939);
and gate_3913(n3941,n3921,n3940);
not gate_3914(n3942,n3941);
and gate_3915(n3943,n30,n3942);
not gate_3916(n3944,n3943);
and gate_3917(n3945,n3899,n3944);
not gate_3918(n3946,n3945);
and gate_3919(n3947,pi1,n3946);
not gate_3920(n3948,n3947);
and gate_3921(n3949,n33,n99);
not gate_3922(n3950,n3949);
and gate_3923(n3951,n1007,n1299);
not gate_3924(n3952,n3951);
and gate_3925(n3953,n3950,n3952);
not gate_3926(n3954,n3953);
and gate_3927(n3955,pi0,n3954);
not gate_3928(n3956,n3955);
and gate_3929(n3957,n132,n1305);
not gate_3930(n3958,n3957);
and gate_3931(n3959,n30,n3958);
not gate_3932(n3960,n3959);
and gate_3933(n3961,n791,n3960);
and gate_3934(n3962,n3956,n3961);
not gate_3935(n3963,n3962);
and gate_3936(n3964,pi4,n3963);
not gate_3937(n3965,n3964);
and gate_3938(n3966,n1693,n2651);
and gate_3939(n3967,n1005,n3966);
and gate_3940(n3968,n38,n3967);
not gate_3941(n3969,n3968);
and gate_3942(n3970,n219,n454);
and gate_3943(n3971,pi0,n3970);
not gate_3944(n3972,n3971);
and gate_3945(n3973,n3969,n3972);
not gate_3946(n3974,n3973);
and gate_3947(n3975,n34,n3974);
not gate_3948(n3976,n3975);
and gate_3949(n3977,n790,n2678);
not gate_3950(n3978,n3977);
and gate_3951(n3979,n3976,n3978);
and gate_3952(n3980,n3965,n3979);
not gate_3953(n3981,n3980);
and gate_3954(n3982,pi2,n3981);
not gate_3955(n3983,n3982);
and gate_3956(n3984,n69,n3421);
not gate_3957(n3985,n3984);
and gate_3958(n3986,n3983,n3985);
not gate_3959(n3987,n3986);
and gate_3960(n3988,n31,n3987);
not gate_3961(n3989,n3988);
and gate_3962(n3990,n821,n2681);
and gate_3963(n3991,n2998,n3990);
not gate_3964(n3992,n3991);
and gate_3965(n3993,n3989,n3992);
and gate_3966(n3994,n3948,n3993);
and gate_3967(n3995,n3862,n3994);
and gate_3968(n3996,n3850,n3995);
not gate_3969(n3997,n3996);
and gate_3970(n3998,pi6,n3997);
not gate_3971(n3999,n3998);
and gate_3972(n4000,n762,n1252);
and gate_3973(n4001,n30,n4000);
not gate_3974(n4002,n4001);
and gate_3975(n4003,n34,n1004);
and gate_3976(n4004,n1243,n4003);
not gate_3977(n4005,n4004);
and gate_3978(n4006,n4002,n4005);
not gate_3979(n4007,n4006);
and gate_3980(n4008,pi3,n4007);
not gate_3981(n4009,n4008);
and gate_3982(n4010,n1215,n1754);
not gate_3983(n4011,n4010);
and gate_3984(n4012,n1184,n1841);
not gate_3985(n4013,n4012);
and gate_3986(n4014,n4011,n4013);
not gate_3987(n4015,n4014);
and gate_3988(n4016,n897,n4015);
not gate_3989(n4017,n4016);
and gate_3990(n4018,n4009,n4017);
and gate_3991(n4019,n37,n1085);
not gate_3992(n4020,n4019);
and gate_3993(n4021,n1186,n4020);
and gate_3994(n4022,n30,n4021);
not gate_3995(n4023,n4022);
and gate_3996(n4024,n30,n1079);
not gate_3997(n4025,n4024);
and gate_3998(n4026,n32,n4025);
not gate_3999(n4027,n4026);
and gate_4000(n4028,n1004,n1184);
not gate_4001(n4029,n4028);
and gate_4002(n4030,n4027,n4029);
and gate_4003(n4031,n4023,n4030);
not gate_4004(n4032,n4031);
and gate_4005(n4033,n38,n4032);
not gate_4006(n4034,n4033);
and gate_4007(n4035,n257,n2093);
not gate_4008(n4036,n4035);
and gate_4009(n4037,n286,n2325);
not gate_4010(n4038,n4037);
and gate_4011(n4039,n1974,n4038);
and gate_4012(n4040,n3085,n4039);
not gate_4013(n4041,n4040);
and gate_4014(n4042,n4036,n4041);
and gate_4015(n4043,n4034,n4042);
not gate_4016(n4044,n4043);
and gate_4017(n4045,pi1,n4044);
not gate_4018(n4046,n4045);
and gate_4019(n4047,pi4,n2746);
not gate_4020(n4048,n4047);
and gate_4021(n4049,n54,n4048);
and gate_4022(n4050,n31,n4049);
not gate_4023(n4051,n4050);
and gate_4024(n4052,n32,n480);
not gate_4025(n4053,n4052);
and gate_4026(n4054,n4051,n4053);
not gate_4027(n4055,n4054);
and gate_4028(n4056,n35,n4055);
not gate_4029(n4057,n4056);
and gate_4030(n4058,n512,n2698);
and gate_4031(n4059,n31,n4058);
not gate_4032(n4060,n4059);
and gate_4033(n4061,n4057,n4060);
not gate_4034(n4062,n4061);
and gate_4035(n4063,pi0,n4062);
not gate_4036(n4064,n4063);
and gate_4037(n4065,n454,n663);
and gate_4038(n4066,n695,n4065);
and gate_4039(n4067,n31,n4066);
not gate_4040(n4068,n4067);
and gate_4041(n4069,n81,n509);
not gate_4042(n4070,n4069);
and gate_4043(n4071,n4068,n4070);
not gate_4044(n4072,n4071);
and gate_4045(n4073,n30,n4072);
not gate_4046(n4074,n4073);
and gate_4047(n4075,n131,n2825);
not gate_4048(n4076,n4075);
and gate_4049(n4077,n4074,n4076);
not gate_4050(n4078,n4077);
and gate_4051(n4079,pi2,n4078);
not gate_4052(n4080,n4079);
and gate_4053(n4081,n4064,n4080);
and gate_4054(n4082,n4046,n4081);
not gate_4055(n4083,n4082);
and gate_4056(n4084,n33,n4083);
not gate_4057(n4085,n4084);
and gate_4058(n4086,n1288,n1327);
not gate_4059(n4087,n4086);
and gate_4060(n4088,n31,n4087);
not gate_4061(n4089,n4088);
and gate_4062(n4090,n563,n2892);
and gate_4063(n4091,n4089,n4090);
not gate_4064(n4092,n4091);
and gate_4065(n4093,pi2,n4092);
not gate_4066(n4094,n4093);
and gate_4067(n4095,n82,n1274);
not gate_4068(n4096,n4095);
and gate_4069(n4097,pi1,n4096);
not gate_4070(n4098,n4097);
and gate_4071(n4099,n1195,n4098);
not gate_4072(n4100,n4099);
and gate_4073(n4101,n32,n4100);
not gate_4074(n4102,n4101);
and gate_4075(n4103,n4094,n4102);
not gate_4076(n4104,n4103);
and gate_4077(n4105,pi5,n4104);
not gate_4078(n4106,n4105);
and gate_4079(n4107,n129,n2870);
not gate_4080(n4108,n4107);
and gate_4081(n4109,n1288,n4108);
not gate_4082(n4110,n4109);
and gate_4083(n4111,pi1,n4110);
not gate_4084(n4112,n4111);
and gate_4085(n4113,n37,n968);
and gate_4086(n4114,n32,n4113);
not gate_4087(n4115,n4114);
and gate_4088(n4116,n35,n3489);
and gate_4089(n4117,n31,n4116);
not gate_4090(n4118,n4117);
and gate_4091(n4119,n4115,n4118);
not gate_4092(n4120,n4119);
and gate_4093(n4121,pi4,n4120);
not gate_4094(n4122,n4121);
and gate_4095(n4123,n4112,n4122);
and gate_4096(n4124,n4106,n4123);
not gate_4097(n4125,n4124);
and gate_4098(n4126,pi0,n4125);
not gate_4099(n4127,n4126);
and gate_4100(n4128,n887,n1365);
not gate_4101(n4129,n4128);
and gate_4102(n4130,n82,n4129);
and gate_4103(n4131,n30,n4130);
not gate_4104(n4132,n4131);
and gate_4105(n4133,pi8,n888);
and gate_4106(n4134,n2826,n4133);
not gate_4107(n4135,n4134);
and gate_4108(n4136,n4132,n4135);
not gate_4109(n4137,n4136);
and gate_4110(n4138,n35,n4137);
not gate_4111(n4139,n4138);
and gate_4112(n4140,n560,n1586);
not gate_4113(n4141,n4140);
and gate_4114(n4142,n4139,n4141);
not gate_4115(n4143,n4142);
and gate_4116(n4144,pi2,n4143);
not gate_4117(n4145,n4144);
and gate_4118(n4146,n4127,n4145);
not gate_4119(n4147,n4146);
and gate_4120(n4148,pi3,n4147);
not gate_4121(n4149,n4148);
and gate_4122(n4150,n32,n694);
not gate_4123(n4151,n4150);
and gate_4124(n4152,n639,n4150);
not gate_4125(n4153,n4152);
and gate_4126(n4154,n4108,n4153);
not gate_4127(n4155,n4154);
and gate_4128(n4156,n31,n4155);
not gate_4129(n4157,n4156);
and gate_4130(n4158,n1347,n2857);
not gate_4131(n4159,n4158);
and gate_4132(n4160,n4157,n4159);
not gate_4133(n4161,n4160);
and gate_4134(n4162,pi0,n4161);
not gate_4135(n4163,n4162);
and gate_4136(n4164,n4149,n4163);
and gate_4137(n4165,n4085,n4164);
and gate_4138(n4166,n4018,n4165);
not gate_4139(n4167,n4166);
and gate_4140(n4168,n36,n4167);
not gate_4141(n4169,n4168);
and gate_4142(n4170,n1692,n2857);
not gate_4143(n4171,n4170);
and gate_4144(n4172,pi0,n1128);
not gate_4145(n4173,n4172);
and gate_4146(n4174,n30,n1004);
not gate_4147(n4175,n4174);
and gate_4148(n4176,n4173,n4175);
not gate_4149(n4177,n4176);
and gate_4150(n4178,n1299,n4177);
not gate_4151(n4179,n4178);
and gate_4152(n4180,n4171,n4179);
not gate_4153(n4181,n4180);
and gate_4154(n4182,n32,n4181);
not gate_4155(n4183,n4182);
and gate_4156(n4184,n39,n1577);
not gate_4157(n4185,n4184);
and gate_4158(n4186,n4183,n4185);
not gate_4159(n4187,n4186);
and gate_4160(n4188,pi1,n4187);
not gate_4161(n4189,n4188);
and gate_4162(n4190,n801,n2857);
not gate_4163(n4191,n4190);
and gate_4164(n4192,n4189,n4191);
not gate_4165(n4193,n4192);
and gate_4166(n4194,n34,n4193);
not gate_4167(n4195,n4194);
and gate_4168(n4196,n4169,n4195);
and gate_4169(n4197,n3999,n4196);
not gate_4170(po10,n4197);
and gate_4171(n4199,n1259,n1430);
not gate_4172(n4200,n4199);
and gate_4173(n4201,n563,n1431);
not gate_4174(n4202,n4201);
and gate_4175(n4203,pi0,n4202);
not gate_4176(n4204,n4203);
and gate_4177(n4205,n43,n1552);
not gate_4178(n4206,n4205);
and gate_4179(n4207,n4204,n4206);
not gate_4180(n4208,n4207);
and gate_4181(n4209,n1145,n4208);
not gate_4182(n4210,n4209);
and gate_4183(n4211,n4200,n4210);
not gate_4184(n4212,n4211);
and gate_4185(n4213,pi6,n4212);
not gate_4186(n4214,n4213);
and gate_4187(n4215,n39,n422);
not gate_4188(n4216,n4215);
and gate_4189(n4217,n1259,n4215);
not gate_4190(n4218,n4217);
and gate_4191(n4219,n4214,n4218);
not gate_4192(n4220,n4219);
and gate_4193(n4221,n1254,n4220);
not gate_4194(n4222,n4221);
and gate_4195(n4223,n223,n1203);
and gate_4196(n4224,n150,n4223);
and gate_4197(n4225,n30,n4224);
not gate_4198(n4226,n4225);
and gate_4199(n4227,pi0,n953);
and gate_4200(n4228,n998,n4227);
not gate_4201(n4229,n4228);
and gate_4202(n4230,n4226,n4229);
not gate_4203(n4231,n4230);
and gate_4204(n4232,pi2,n4231);
not gate_4205(n4233,n4232);
and gate_4206(n4234,n30,n1145);
and gate_4207(n4235,n179,n519);
and gate_4208(n4236,n4234,n4235);
not gate_4209(n4237,n4236);
and gate_4210(n4238,n4233,n4237);
not gate_4211(n4239,n4238);
and gate_4212(n4240,n639,n4239);
not gate_4213(n4241,n4240);
and gate_4214(n4242,n291,n642);
not gate_4215(n4243,n4242);
and gate_4216(n4244,n644,n897);
not gate_4217(n4245,n4244);
and gate_4218(n4246,n4243,n4245);
not gate_4219(n4247,n4246);
and gate_4220(n4248,pi0,n4247);
not gate_4221(n4249,n4248);
and gate_4222(n4250,pi4,n181);
and gate_4223(n4251,n3741,n4250);
not gate_4224(n4252,n4251);
and gate_4225(n4253,n4249,n4252);
not gate_4226(n4254,n4253);
and gate_4227(n4255,n35,n4254);
not gate_4228(n4256,n4255);
and gate_4229(n4257,n179,n1363);
not gate_4230(n4258,n4257);
and gate_4231(n4259,n181,n435);
not gate_4232(n4260,n4259);
and gate_4233(n4261,n4258,n4260);
not gate_4234(n4262,n4261);
and gate_4235(n4263,n116,n4262);
not gate_4236(n4264,n4263);
and gate_4237(n4265,n4256,n4264);
not gate_4238(n4266,n4265);
and gate_4239(n4267,pi2,n4266);
not gate_4240(n4268,n4267);
and gate_4241(n4269,n998,n2555);
not gate_4242(n4270,n4269);
and gate_4243(n4271,n1008,n2562);
not gate_4244(n4272,n4271);
and gate_4245(n4273,n4270,n4272);
not gate_4246(n4274,n4273);
and gate_4247(n4275,n817,n4274);
not gate_4248(n4276,n4275);
and gate_4249(n4277,n4268,n4276);
and gate_4250(n4278,n32,n1078);
not gate_4251(n4279,n4278);
and gate_4252(n4280,n1453,n4279);
not gate_4253(n4281,n4280);
and gate_4254(n4282,n34,n663);
not gate_4255(n4283,n4282);
and gate_4256(n4284,pi1,n4283);
not gate_4257(n4285,n4284);
and gate_4258(n4286,n785,n4285);
not gate_4259(n4287,n4286);
and gate_4260(n4288,n1049,n4287);
and gate_4261(n4289,n4281,n4288);
not gate_4262(n4290,n4289);
and gate_4263(n4291,n181,n1577);
not gate_4264(n4292,n4291);
and gate_4265(n4293,n1176,n3320);
not gate_4266(n4294,n4293);
and gate_4267(n4295,n4292,n4294);
not gate_4268(n4296,n4295);
and gate_4269(n4297,n31,n451);
not gate_4270(n4298,n4297);
and gate_4271(n4299,pi1,n636);
not gate_4272(n4300,n4299);
and gate_4273(n4301,n4298,n4300);
not gate_4274(n4302,n4301);
and gate_4275(n4303,n4296,n4302);
not gate_4276(n4304,n4303);
and gate_4277(n4305,n97,n1577);
not gate_4278(n4306,n4305);
and gate_4279(n4307,n117,n1100);
not gate_4280(n4308,n4307);
and gate_4281(n4309,n4306,n4308);
not gate_4282(n4310,n4309);
and gate_4283(n4311,pi1,n4310);
not gate_4284(n4312,n4311);
and gate_4285(n4313,n1854,n3438);
and gate_4286(n4314,n31,n4313);
not gate_4287(n4315,n4314);
and gate_4288(n4316,n4312,n4315);
not gate_4289(n4317,n4316);
and gate_4290(n4318,pi4,n4317);
not gate_4291(n4319,n4318);
and gate_4292(n4320,n32,n3151);
not gate_4293(n4321,n4320);
and gate_4294(n4322,pi2,n181);
not gate_4295(n4323,n4322);
and gate_4296(n4324,n4321,n4323);
not gate_4297(n4325,n4324);
and gate_4298(n4326,n35,n4325);
not gate_4299(n4327,n4326);
and gate_4300(n4328,n43,n1918);
not gate_4301(n4329,n4328);
and gate_4302(n4330,n4327,n4329);
not gate_4303(n4331,n4330);
and gate_4304(n4332,n435,n4331);
not gate_4305(n4333,n4332);
and gate_4306(n4334,n4319,n4333);
and gate_4307(n4335,n4304,n4334);
and gate_4308(n4336,n4290,n4335);
not gate_4309(n4337,n4336);
and gate_4310(n4338,pi0,n4337);
not gate_4311(n4339,n4338);
and gate_4312(n4340,pi4,n259);
and gate_4313(n4341,n853,n4340);
not gate_4314(n4342,n4341);
and gate_4315(n4343,n436,n4342);
not gate_4316(n4344,n4343);
and gate_4317(n4345,n35,n4344);
not gate_4318(n4346,n4345);
and gate_4319(n4347,n560,n1363);
not gate_4320(n4348,n4347);
and gate_4321(n4349,n4346,n4348);
not gate_4322(n4350,n4349);
and gate_4323(n4351,pi6,n4350);
not gate_4324(n4352,n4351);
and gate_4325(n4353,n175,n4134);
not gate_4326(n4354,n4353);
and gate_4327(n4355,n4352,n4354);
not gate_4328(n4356,n4355);
and gate_4329(n4357,pi2,n4356);
not gate_4330(n4358,n4357);
and gate_4331(n4359,n790,n1145);
not gate_4332(n4360,n4359);
and gate_4333(n4361,pi1,n4360);
not gate_4334(n4362,n4361);
and gate_4335(n4363,n34,n4362);
not gate_4336(n4364,n4363);
and gate_4337(n4365,n270,n707);
not gate_4338(n4366,n4365);
and gate_4339(n4367,n1347,n4366);
not gate_4340(n4368,n4367);
and gate_4341(n4369,n4364,n4368);
not gate_4342(n4370,n4369);
and gate_4343(n4371,n36,n4370);
not gate_4344(n4372,n4371);
and gate_4345(n4373,n4358,n4372);
not gate_4346(n4374,n4373);
and gate_4347(n4375,n30,n4374);
not gate_4348(n4376,n4375);
and gate_4349(n4377,n31,n1184);
and gate_4350(n4378,n152,n4377);
not gate_4351(n4379,n4378);
and gate_4352(n4380,n4376,n4379);
and gate_4353(n4381,n4339,n4380);
not gate_4354(n4382,n4381);
and gate_4355(n4383,n33,n4382);
not gate_4356(n4384,n4383);
and gate_4357(n4385,n762,n4234);
not gate_4358(n4386,n4385);
and gate_4359(n4387,n2562,n4281);
not gate_4360(n4388,n4387);
and gate_4361(n4389,n4386,n4388);
not gate_4362(n4390,n4389);
and gate_4363(n4391,n2198,n4390);
not gate_4364(n4392,n4391);
and gate_4365(n4393,n37,n456);
not gate_4366(n4394,n4393);
and gate_4367(n4395,n4065,n4394);
and gate_4368(n4396,pi1,n4395);
not gate_4369(n4397,n4396);
and gate_4370(n4398,n1895,n4397);
not gate_4371(n4399,n4398);
and gate_4372(n4400,n32,n4399);
not gate_4373(n4401,n4400);
and gate_4374(n4402,pi2,n460);
not gate_4375(n4403,n4402);
and gate_4376(n4404,n590,n1182);
not gate_4377(n4405,n4404);
and gate_4378(n4406,n4403,n4405);
not gate_4379(n4407,n4406);
and gate_4380(n4408,n852,n4407);
not gate_4381(n4409,n4408);
and gate_4382(n4410,n4401,n4409);
not gate_4383(n4411,n4410);
and gate_4384(n4412,n36,n4411);
not gate_4385(n4413,n4412);
and gate_4386(n4414,n34,n268);
not gate_4387(n4415,n4414);
and gate_4388(n4416,n1431,n4415);
not gate_4389(n4417,n4416);
and gate_4390(n4418,n35,n4417);
not gate_4391(n4419,n4418);
and gate_4392(n4420,n277,n3139);
not gate_4393(n4421,n4420);
and gate_4394(n4422,n4419,n4421);
not gate_4395(n4423,n4422);
and gate_4396(n4424,pi6,n4423);
and gate_4397(n4425,n1137,n4424);
not gate_4398(n4426,n4425);
and gate_4399(n4427,n4413,n4426);
not gate_4400(n4428,n4427);
and gate_4401(n4429,pi0,n4428);
not gate_4402(n4430,n4429);
and gate_4403(n4431,n104,n4283);
and gate_4404(n4432,n32,n4431);
not gate_4405(n4433,n4432);
and gate_4406(n4434,n885,n1286);
not gate_4407(n4435,n4434);
and gate_4408(n4436,n3051,n4435);
not gate_4409(n4437,n4436);
and gate_4410(n4438,n4433,n4437);
not gate_4411(n4439,n4438);
and gate_4412(n4440,n35,n4439);
not gate_4413(n4441,n4440);
and gate_4414(n4442,pi2,n509);
not gate_4415(n4443,n4442);
and gate_4416(n4444,n1183,n4443);
not gate_4417(n4445,n4444);
and gate_4418(n4446,n117,n4445);
not gate_4419(n4447,n4446);
and gate_4420(n4448,n4441,n4447);
not gate_4421(n4449,n4448);
and gate_4422(n4450,n1586,n4449);
not gate_4423(n4451,n4450);
and gate_4424(n4452,n4430,n4451);
and gate_4425(n4453,n4392,n4452);
not gate_4426(n4454,n4453);
and gate_4427(n4455,pi3,n4454);
not gate_4428(n4456,n4455);
and gate_4429(n4457,n299,n1078);
not gate_4430(n4458,n4457);
and gate_4431(n4459,pi1,n4150);
not gate_4432(n4460,n4459);
and gate_4433(n4461,n4458,n4460);
not gate_4434(n4462,n4461);
and gate_4435(n4463,n3677,n4462);
and gate_4436(n4464,pi0,n4463);
not gate_4437(n4465,n4464);
and gate_4438(n4466,n30,n1241);
not gate_4439(n4467,n4466);
and gate_4440(n4468,n4465,n4467);
and gate_4441(n4469,n4456,n4468);
and gate_4442(n4470,n4384,n4469);
and gate_4443(n4471,n4277,n4470);
and gate_4444(n4472,n4241,n4471);
and gate_4445(n4473,n4222,n4472);
not gate_4446(po11,n4473);
and gate_4447(n4475,pi2,n4414);
not gate_4448(n4476,n4475);
and gate_4449(n4477,n43,n1182);
not gate_4450(n4478,n4477);
and gate_4451(n4479,n4476,n4478);
not gate_4452(n4480,n4479);
and gate_4453(n4481,n178,n4480);
not gate_4454(n4482,n4481);
and gate_4455(n4483,pi2,n277);
and gate_4456(n4484,n117,n4483);
not gate_4457(n4485,n4484);
and gate_4458(n4486,n39,n626);
not gate_4459(n4487,n4486);
and gate_4460(n4488,n43,n784);
not gate_4461(n4489,n4488);
and gate_4462(n4490,n4487,n4489);
not gate_4463(n4491,n4490);
and gate_4464(n4492,n1100,n4491);
not gate_4465(n4493,n4492);
and gate_4466(n4494,n4485,n4493);
and gate_4467(n4495,n4482,n4494);
not gate_4468(n4496,n4495);
and gate_4469(n4497,n31,n4496);
not gate_4470(n4498,n4497);
and gate_4471(n4499,n179,n1100);
not gate_4472(n4500,n4499);
and gate_4473(n4501,n4292,n4500);
and gate_4474(n4502,n1186,n3445);
and gate_4475(n4503,n191,n4502);
not gate_4476(n4504,n4503);
and gate_4477(n4505,n4501,n4504);
not gate_4478(n4506,n4505);
and gate_4479(n4507,pi8,n4506);
not gate_4480(n4508,n4507);
and gate_4481(n4509,n1101,n3052);
not gate_4482(n4510,n4509);
and gate_4483(n4511,n1006,n4510);
and gate_4484(n4512,n38,n4511);
not gate_4485(n4513,n4512);
and gate_4486(n4514,n104,n1577);
not gate_4487(n4515,n4514);
and gate_4488(n4516,n4513,n4515);
not gate_4489(n4517,n4516);
and gate_4490(n4518,pi4,n4517);
not gate_4491(n4519,n4518);
and gate_4492(n4520,n34,n4307);
not gate_4493(n4521,n4520);
and gate_4494(n4522,n4519,n4521);
and gate_4495(n4523,n4508,n4522);
not gate_4496(n4524,n4523);
and gate_4497(n4525,pi1,n4524);
not gate_4498(n4526,n4525);
and gate_4499(n4527,n4498,n4526);
not gate_4500(n4528,n4527);
and gate_4501(n4529,pi3,n4528);
not gate_4502(n4530,n4529);
and gate_4503(n4531,pi4,n1078);
not gate_4504(n4532,n4531);
and gate_4505(n4533,n4151,n4532);
not gate_4506(n4534,n4533);
and gate_4507(n4535,n1183,n4534);
and gate_4508(n4536,pi1,n4535);
not gate_4509(n4537,n4536);
and gate_4510(n4538,n299,n762);
not gate_4511(n4539,n4538);
and gate_4512(n4540,n4537,n4539);
not gate_4513(n4541,n4540);
and gate_4514(n4542,pi6,n4541);
not gate_4515(n4543,n4542);
and gate_4516(n4544,n1614,n2516);
not gate_4517(n4545,n4544);
and gate_4518(n4546,n4543,n4545);
and gate_4519(n4547,n1181,n4302);
not gate_4520(n4548,n4547);
and gate_4521(n4549,pi2,n886);
not gate_4522(n4550,n4549);
and gate_4523(n4551,n563,n4550);
not gate_4524(n4552,n4551);
and gate_4525(n4553,pi1,n4552);
not gate_4526(n4554,n4553);
and gate_4527(n4555,n4548,n4554);
not gate_4528(n4556,n4555);
and gate_4529(n4557,n36,n4556);
not gate_4530(n4558,n4557);
and gate_4531(n4559,n1137,n3421);
not gate_4532(n4560,n4559);
and gate_4533(n4561,n40,n1431);
not gate_4534(n4562,n4561);
and gate_4535(n4563,n1241,n4562);
not gate_4536(n4564,n4563);
and gate_4537(n4565,n4560,n4564);
not gate_4538(n4566,n4565);
and gate_4539(n4567,pi6,n4566);
not gate_4540(n4568,n4567);
and gate_4541(n4569,n4558,n4568);
not gate_4542(n4570,n4569);
and gate_4543(n4571,pi5,n4570);
not gate_4544(n4572,n4571);
and gate_4545(n4573,n31,n1178);
not gate_4546(n4574,n4573);
and gate_4547(n4575,n268,n1145);
and gate_4548(n4576,n36,n4575);
not gate_4549(n4577,n4576);
and gate_4550(n4578,n4574,n4577);
not gate_4551(n4579,n4578);
and gate_4552(n4580,n608,n4579);
not gate_4553(n4581,n4580);
and gate_4554(n4582,n4572,n4581);
and gate_4555(n4583,n4546,n4582);
not gate_4556(n4584,n4583);
and gate_4557(n4585,n33,n4584);
not gate_4558(n4586,n4585);
and gate_4559(n4587,n4530,n4586);
not gate_4560(n4588,n4587);
and gate_4561(n4589,pi0,n4588);
not gate_4562(n4590,n4589);
and gate_4563(n4591,n435,n1167);
not gate_4564(n4592,n4591);
and gate_4565(n4593,pi1,n178);
not gate_4566(n4594,n4593);
and gate_4567(n4595,n31,n150);
not gate_4568(n4596,n4595);
and gate_4569(n4597,n4594,n4596);
not gate_4570(n4598,n4597);
and gate_4571(n4599,n257,n4598);
not gate_4572(n4600,n4599);
and gate_4573(n4601,n4592,n4600);
not gate_4574(n4602,n4601);
and gate_4575(n4603,pi2,n4602);
not gate_4576(n4604,n4603);
and gate_4577(n4605,n32,n2042);
and gate_4578(n4606,n2891,n4605);
not gate_4579(n4607,n4606);
and gate_4580(n4608,n4604,n4607);
and gate_4581(n4609,n43,n424);
not gate_4582(n4610,n4609);
and gate_4583(n4611,n4216,n4610);
not gate_4584(n4612,n4611);
and gate_4585(n4613,n31,n4612);
not gate_4586(n4614,n4613);
and gate_4587(n4615,n587,n869);
not gate_4588(n4616,n4615);
and gate_4589(n4617,n4614,n4616);
not gate_4590(n4618,n4617);
and gate_4591(n4619,n1577,n4618);
not gate_4592(n4620,n4619);
and gate_4593(n4621,n42,n44);
not gate_4594(n4622,n4621);
and gate_4595(n4623,n608,n4622);
and gate_4596(n4624,n1145,n4623);
not gate_4597(n4625,n4624);
and gate_4598(n4626,n4620,n4625);
and gate_4599(n4627,n4608,n4626);
not gate_4600(n4628,n4627);
and gate_4601(n4629,pi3,n4628);
not gate_4602(n4630,n4629);
and gate_4603(n4631,pi2,n1874);
not gate_4604(n4632,n4631);
and gate_4605(n4633,n1223,n4632);
not gate_4606(n4634,n4633);
and gate_4607(n4635,n37,n4634);
not gate_4608(n4636,n4635);
and gate_4609(n4637,n1176,n2043);
not gate_4610(n4638,n4637);
and gate_4611(n4639,n4636,n4638);
not gate_4612(n4640,n4639);
and gate_4613(n4641,n34,n4640);
not gate_4614(n4642,n4641);
and gate_4615(n4643,pi2,n271);
not gate_4616(n4644,n4643);
and gate_4617(n4645,n4642,n4644);
not gate_4618(n4646,n4645);
and gate_4619(n4647,pi1,n4646);
not gate_4620(n4648,n4647);
and gate_4621(n4649,n425,n1431);
not gate_4622(n4650,n4649);
and gate_4623(n4651,pi5,n3422);
not gate_4624(n4652,n4651);
and gate_4625(n4653,n4650,n4652);
and gate_4626(n4654,pi2,n4653);
not gate_4627(n4655,n4654);
and gate_4628(n4656,pi4,n130);
not gate_4629(n4657,n4656);
and gate_4630(n4658,n36,n4657);
not gate_4631(n4659,n4658);
and gate_4632(n4660,n4655,n4659);
not gate_4633(n4661,n4660);
and gate_4634(n4662,n31,n4661);
not gate_4635(n4663,n4662);
and gate_4636(n4664,n617,n4442);
not gate_4637(n4665,n4664);
and gate_4638(n4666,n4663,n4665);
and gate_4639(n4667,n4648,n4666);
not gate_4640(n4668,n4667);
and gate_4641(n4669,n33,n4668);
not gate_4642(n4670,n4669);
and gate_4643(n4671,n1242,n4670);
and gate_4644(n4672,n4630,n4671);
not gate_4645(n4673,n4672);
and gate_4646(n4674,n30,n4673);
not gate_4647(n4675,n4674);
and gate_4648(n4676,n4590,n4675);
not gate_4649(po12,n4676);
and gate_4650(n4678,n596,n1192);
not gate_4651(n4679,n4678);
and gate_4652(n4680,n1154,n1634);
not gate_4653(n4681,n4680);
and gate_4654(n4682,n4679,n4681);
not gate_4655(n4683,n4682);
and gate_4656(n4684,n31,n4683);
not gate_4657(n4685,n4684);
and gate_4658(n4686,n1490,n1703);
and gate_4659(n4687,n1137,n4686);
not gate_4660(n4688,n4687);
and gate_4661(n4689,n4685,n4688);
not gate_4662(n4690,n4689);
and gate_4663(n4691,pi0,n4690);
not gate_4664(n4692,n4691);
and gate_4665(n4693,n819,n2834);
not gate_4666(n4694,n4693);
and gate_4667(n4695,n114,n1145);
not gate_4668(n4696,n4695);
and gate_4669(n4697,n4694,n4696);
not gate_4670(n4698,n4697);
and gate_4671(n4699,n1552,n4698);
not gate_4672(n4700,n4699);
and gate_4673(n4701,n4692,n4700);
not gate_4674(n4702,n4701);
and gate_4675(n4703,n37,n4702);
not gate_4676(n4704,n4703);
and gate_4677(n4705,n926,n4234);
not gate_4678(n4706,n4705);
and gate_4679(n4707,n457,n1154);
not gate_4680(n4708,n4707);
and gate_4681(n4709,n1192,n2818);
not gate_4682(n4710,n4709);
and gate_4683(n4711,n4708,n4710);
not gate_4684(n4712,n4711);
and gate_4685(n4713,n2243,n4712);
not gate_4686(n4714,n4713);
and gate_4687(n4715,n4706,n4714);
not gate_4688(n4716,n4715);
and gate_4689(n4717,pi7,n4716);
not gate_4690(n4718,n4717);
and gate_4691(n4719,n4704,n4718);
and gate_4692(n4720,n30,n200);
not gate_4693(n4721,n4720);
and gate_4694(n4722,pi0,n202);
not gate_4695(n4723,n4722);
and gate_4696(n4724,n4721,n4723);
not gate_4697(n4725,n4724);
and gate_4698(n4726,n4302,n4725);
not gate_4699(n4727,n4726);
and gate_4700(n4728,n313,n3421);
not gate_4701(n4729,n4728);
and gate_4702(n4730,n1326,n2395);
not gate_4703(n4731,n4730);
and gate_4704(n4732,n4729,n4731);
not gate_4705(n4733,n4732);
and gate_4706(n4734,pi3,n4733);
not gate_4707(n4735,n4734);
and gate_4708(n4736,n4727,n4735);
not gate_4709(n4737,n4736);
and gate_4710(n4738,pi2,n4737);
not gate_4711(n4739,n4738);
and gate_4712(n4740,n43,n142);
and gate_4713(n4741,n4234,n4740);
not gate_4714(n4742,n4741);
and gate_4715(n4743,n4739,n4742);
not gate_4716(n4744,n4743);
and gate_4717(n4745,n178,n4744);
not gate_4718(n4746,n4745);
and gate_4719(n4747,n81,n114);
not gate_4720(n4748,n4747);
and gate_4721(n4749,n520,n4748);
not gate_4722(n4750,n4749);
and gate_4723(n4751,n31,n4750);
not gate_4724(n4752,n4751);
and gate_4725(n4753,n62,n217);
and gate_4726(n4754,pi1,n4753);
not gate_4727(n4755,n4754);
and gate_4728(n4756,n4752,n4755);
not gate_4729(n4757,n4756);
and gate_4730(n4758,pi2,n4757);
not gate_4731(n4759,n4758);
and gate_4732(n4760,pi1,n817);
not gate_4733(n4761,n4760);
and gate_4734(n4762,n708,n4760);
not gate_4735(n4763,n4762);
and gate_4736(n4764,n4759,n4763);
not gate_4737(n4765,n4764);
and gate_4738(n4766,n30,n4765);
not gate_4739(n4767,n4766);
and gate_4740(n4768,n114,n260);
not gate_4741(n4769,n4768);
and gate_4742(n4770,n519,n3139);
not gate_4743(n4771,n4770);
and gate_4744(n4772,n4769,n4771);
not gate_4745(n4773,n4772);
and gate_4746(n4774,n32,n4773);
not gate_4747(n4775,n4774);
and gate_4748(n4776,n790,n819);
not gate_4749(n4777,n4776);
and gate_4750(n4778,n4775,n4777);
not gate_4751(n4779,n4778);
and gate_4752(n4780,n2395,n4779);
not gate_4753(n4781,n4780);
and gate_4754(n4782,n4767,n4781);
not gate_4755(n4783,n4782);
and gate_4756(n4784,n34,n4783);
not gate_4757(n4785,n4784);
and gate_4758(n4786,n1007,n1253);
and gate_4759(n4787,n1243,n4786);
not gate_4760(n4788,n4787);
and gate_4761(n4789,n1004,n1137);
and gate_4762(n4790,n2678,n4789);
not gate_4763(n4791,n4790);
and gate_4764(n4792,n4788,n4791);
and gate_4765(n4793,n1299,n2135);
and gate_4766(n4794,pi0,n4793);
not gate_4767(n4795,n4794);
and gate_4768(n4796,n313,n3885);
not gate_4769(n4797,n4796);
and gate_4770(n4798,n4795,n4797);
not gate_4771(n4799,n4798);
and gate_4772(n4800,n35,n4799);
not gate_4773(n4801,n4800);
and gate_4774(n4802,n3822,n4234);
not gate_4775(n4803,n4802);
and gate_4776(n4804,n4801,n4803);
not gate_4777(n4805,n4804);
and gate_4778(n4806,n37,n4805);
not gate_4779(n4807,n4806);
and gate_4780(n4808,n39,n217);
and gate_4781(n4809,n1665,n4808);
not gate_4782(n4810,n4809);
and gate_4783(n4811,n4807,n4810);
and gate_4784(n4812,n4792,n4811);
not gate_4785(n4813,n4812);
and gate_4786(n4814,pi4,n4813);
not gate_4787(n4815,n4814);
and gate_4788(n4816,n4785,n4815);
not gate_4789(n4817,n4816);
and gate_4790(n4818,pi6,n4817);
not gate_4791(n4819,n4818);
and gate_4792(n4820,n1025,n1145);
not gate_4793(n4821,n4820);
and gate_4794(n4822,n345,n4573);
not gate_4795(n4823,n4822);
and gate_4796(n4824,n4821,n4823);
not gate_4797(n4825,n4824);
and gate_4798(n4826,n35,n4825);
not gate_4799(n4827,n4826);
and gate_4800(n4828,n4460,n4827);
not gate_4801(n4829,n4828);
and gate_4802(n4830,n34,n4829);
not gate_4803(n4831,n4830);
and gate_4804(n4832,n39,n980);
not gate_4805(n4833,n4832);
and gate_4806(n4834,n43,n239);
not gate_4807(n4835,n4834);
and gate_4808(n4836,n4833,n4835);
not gate_4809(n4837,n4836);
and gate_4810(n4838,n1182,n4837);
not gate_4811(n4839,n4838);
and gate_4812(n4840,n4831,n4839);
not gate_4813(n4841,n4840);
and gate_4814(n4842,pi0,n4841);
not gate_4815(n4843,n4842);
and gate_4816(n4844,n43,n2870);
not gate_4817(n4845,n4844);
and gate_4818(n4846,pi4,n4845);
not gate_4819(n4847,n4846);
and gate_4820(n4848,n31,n4847);
not gate_4821(n4849,n4848);
and gate_4822(n4850,pi2,n1326);
not gate_4823(n4851,n4850);
and gate_4824(n4852,n3416,n4851);
not gate_4825(n4853,n4852);
and gate_4826(n4854,pi1,n4853);
not gate_4827(n4855,n4854);
and gate_4828(n4856,n4849,n4855);
not gate_4829(n4857,n4856);
and gate_4830(n4858,n33,n4857);
not gate_4831(n4859,n4858);
and gate_4832(n4860,n43,n907);
not gate_4833(n4861,n4860);
and gate_4834(n4862,n2870,n3139);
not gate_4835(n4863,n4862);
and gate_4836(n4864,n4861,n4863);
not gate_4837(n4865,n4864);
and gate_4838(n4866,n953,n4865);
not gate_4839(n4867,n4866);
and gate_4840(n4868,n4859,n4867);
not gate_4841(n4869,n4868);
and gate_4842(n4870,n2878,n4869);
not gate_4843(n4871,n4870);
and gate_4844(n4872,n4843,n4871);
not gate_4845(n4873,n4872);
and gate_4846(n4874,n36,n4873);
not gate_4847(n4875,n4874);
and gate_4848(n4876,n4467,n4875);
and gate_4849(n4877,n4819,n4876);
and gate_4850(n4878,n4746,n4877);
and gate_4851(n4879,n4719,n4878);
not gate_4852(po13,n4879);
and gate_4853(n4881,pi2,n636);
not gate_4854(n4882,n4881);
and gate_4855(n4883,n1183,n4882);
not gate_4856(n4884,n4883);
and gate_4857(n4885,pi1,n4884);
not gate_4858(n4886,n4885);
and gate_4859(n4887,n299,n451);
not gate_4860(n4888,n4887);
and gate_4861(n4889,n4886,n4888);
not gate_4862(n4890,n4889);
and gate_4863(n4891,pi6,n4890);
not gate_4864(n4892,n4891);
and gate_4865(n4893,n544,n1145);
not gate_4866(n4894,n4893);
and gate_4867(n4895,n4892,n4894);
not gate_4868(n4896,n4895);
and gate_4869(n4897,n4725,n4896);
not gate_4870(n4898,n4897);
and gate_4871(n4899,n345,n1178);
and gate_4872(n4900,pi0,n4899);
not gate_4873(n4901,n4900);
and gate_4874(n4902,n821,n1489);
and gate_4875(n4903,n2649,n4902);
not gate_4876(n4904,n4903);
and gate_4877(n4905,n4901,n4904);
not gate_4878(n4906,n4905);
and gate_4879(n4907,n36,n4906);
not gate_4880(n4908,n4907);
and gate_4881(n4909,n837,n1192);
and gate_4882(n4910,pi0,n4909);
not gate_4883(n4911,n4910);
and gate_4884(n4912,n4908,n4911);
not gate_4885(n4913,n4912);
and gate_4886(n4914,pi1,n4913);
not gate_4887(n4915,n4914);
and gate_4888(n4916,pi0,n2711);
not gate_4889(n4917,n4916);
and gate_4890(n4918,n1301,n2579);
not gate_4891(n4919,n4918);
and gate_4892(n4920,n4917,n4919);
not gate_4893(n4921,n4920);
and gate_4894(n4922,pi6,n4921);
and gate_4895(n4923,n31,n4922);
not gate_4896(n4924,n4923);
and gate_4897(n4925,n4915,n4924);
and gate_4898(n4926,n617,n869);
not gate_4899(n4927,n4926);
and gate_4900(n4928,n117,n2825);
not gate_4901(n4929,n4928);
and gate_4902(n4930,n4927,n4929);
not gate_4903(n4931,n4930);
and gate_4904(n4932,pi2,n4931);
not gate_4905(n4933,n4932);
and gate_4906(n4934,pi4,n82);
not gate_4907(n4935,n4934);
and gate_4908(n4936,n31,n4935);
not gate_4909(n4937,n4936);
and gate_4910(n4938,n1145,n1326);
not gate_4911(n4939,n4938);
and gate_4912(n4940,n4937,n4939);
not gate_4913(n4941,n4940);
and gate_4914(n4942,n36,n4941);
not gate_4915(n4943,n4942);
and gate_4916(n4944,pi1,n3436);
not gate_4917(n4945,n4944);
and gate_4918(n4946,n3421,n4945);
not gate_4919(n4947,n4946);
and gate_4920(n4948,n4943,n4947);
and gate_4921(n4949,n4933,n4948);
not gate_4922(n4950,n4949);
and gate_4923(n4951,n30,n4950);
not gate_4924(n4952,n4951);
and gate_4925(n4953,n452,n1049);
and gate_4926(n4954,n31,n423);
not gate_4927(n4955,n4954);
and gate_4928(n4956,n4953,n4955);
and gate_4929(n4957,pi7,n4956);
not gate_4930(n4958,n4957);
and gate_4931(n4959,n435,n882);
not gate_4932(n4960,n4959);
and gate_4933(n4961,n4958,n4960);
not gate_4934(n4962,n4961);
and gate_4935(n4963,n32,n4962);
not gate_4936(n4964,n4963);
and gate_4937(n4965,n31,n2870);
not gate_4938(n4966,n4965);
and gate_4939(n4967,n630,n4965);
not gate_4940(n4968,n4967);
and gate_4941(n4969,n4964,n4968);
not gate_4942(n4970,n4969);
and gate_4943(n4971,pi0,n4970);
not gate_4944(n4972,n4971);
and gate_4945(n4973,n4952,n4972);
not gate_4946(n4974,n4973);
and gate_4947(n4975,n33,n4974);
not gate_4948(n4976,n4975);
and gate_4949(n4977,pi2,n104);
not gate_4950(n4978,n4977);
and gate_4951(n4979,n66,n4978);
not gate_4952(n4980,n4979);
and gate_4953(n4981,pi4,n4980);
not gate_4954(n4982,n4981);
and gate_4955(n4983,n3438,n4414);
not gate_4956(n4984,n4983);
and gate_4957(n4985,n4982,n4984);
not gate_4958(n4986,n4985);
and gate_4959(n4987,pi3,n4986);
not gate_4960(n4988,n4987);
and gate_4961(n4989,n617,n2870);
not gate_4962(n4990,n4989);
and gate_4963(n4991,n4988,n4990);
not gate_4964(n4992,n4991);
and gate_4965(n4993,n31,n4992);
not gate_4966(n4994,n4993);
and gate_4967(n4995,n53,n424);
and gate_4968(n4996,n4760,n4995);
not gate_4969(n4997,n4996);
and gate_4970(n4998,n4994,n4997);
not gate_4971(n4999,n4998);
and gate_4972(n5000,pi0,n4999);
not gate_4973(n5001,n5000);
and gate_4974(n5002,n313,n1192);
and gate_4975(n5003,n4215,n5002);
not gate_4976(n5004,n5003);
and gate_4977(n5005,n5001,n5004);
and gate_4978(n5006,n4976,n5005);
and gate_4979(n5007,n4925,n5006);
and gate_4980(n5008,n4898,n5007);
not gate_4981(n5009,n5008);
and gate_4982(n5010,n35,n5009);
not gate_4983(n5011,n5010);
and gate_4984(n5012,pi6,n2708);
not gate_4985(n5013,n5012);
and gate_4986(n5014,n1919,n5013);
not gate_4987(n5015,n5014);
and gate_4988(n5016,pi4,n5015);
not gate_4989(n5017,n5016);
and gate_4990(n5018,n1184,n2198);
not gate_4991(n5019,n5018);
and gate_4992(n5020,n5017,n5019);
not gate_4993(n5021,n5020);
and gate_4994(n5022,n37,n5021);
not gate_4995(n5023,n5022);
and gate_4996(n5024,n2488,n3678);
not gate_4997(n5025,n5024);
and gate_4998(n5026,n2698,n5025);
not gate_4999(n5027,n5026);
and gate_5000(n5028,n5023,n5027);
not gate_5001(n5029,n5028);
and gate_5002(n5030,n33,n5029);
not gate_5003(n5031,n5030);
and gate_5004(n5032,pi4,n2198);
not gate_5005(n5033,n5032);
and gate_5006(n5034,n785,n5033);
not gate_5007(n5035,n5034);
and gate_5008(n5036,n32,n5035);
not gate_5009(n5037,n5036);
and gate_5010(n5038,n332,n1184);
not gate_5011(n5039,n5038);
and gate_5012(n5040,n5037,n5039);
not gate_5013(n5041,n5040);
and gate_5014(n5042,n221,n5041);
not gate_5015(n5043,n5042);
and gate_5016(n5044,n5031,n5043);
not gate_5017(n5045,n5044);
and gate_5018(n5046,n30,n5045);
not gate_5019(n5047,n5046);
and gate_5020(n5048,n104,n206);
not gate_5021(n5049,n5048);
and gate_5022(n5050,n192,n617);
not gate_5023(n5051,n5050);
and gate_5024(n5052,n5049,n5051);
not gate_5025(n5053,n5052);
and gate_5026(n5054,pi2,n5053);
not gate_5027(n5055,n5054);
and gate_5028(n5056,n33,n666);
not gate_5029(n5057,n5056);
and gate_5030(n5058,n37,n345);
not gate_5031(n5059,n5058);
and gate_5032(n5060,n36,n749);
and gate_5033(n5061,n5059,n5060);
not gate_5034(n5062,n5061);
and gate_5035(n5063,n5057,n5062);
not gate_5036(n5064,n5063);
and gate_5037(n5065,pi4,n5064);
not gate_5038(n5066,n5065);
and gate_5039(n5067,n42,n4610);
not gate_5040(n5068,n5067);
and gate_5041(n5069,pi3,n5068);
not gate_5042(n5070,n5069);
and gate_5043(n5071,n5066,n5070);
not gate_5044(n5072,n5071);
and gate_5045(n5073,n32,n5072);
not gate_5046(n5074,n5073);
and gate_5047(n5075,n5055,n5074);
not gate_5048(n5076,n5075);
and gate_5049(n5077,pi0,n5076);
not gate_5050(n5078,n5077);
and gate_5051(n5079,n5047,n5078);
not gate_5052(n5080,n5079);
and gate_5053(n5081,pi1,n5080);
not gate_5054(n5082,n5081);
and gate_5055(n5083,n33,n48);
not gate_5056(n5084,n5083);
and gate_5057(n5085,n53,n225);
not gate_5058(n5086,n5085);
and gate_5059(n5087,n5084,n5086);
not gate_5060(n5088,n5087);
and gate_5061(n5089,pi4,n5088);
not gate_5062(n5090,n5089);
and gate_5063(n5091,n192,n3076);
not gate_5064(n5092,n5091);
and gate_5065(n5093,n5090,n5092);
not gate_5066(n5094,n5093);
and gate_5067(n5095,n30,n5094);
not gate_5068(n5096,n5095);
and gate_5069(n5097,n1265,n2258);
not gate_5070(n5098,n5097);
and gate_5071(n5099,pi3,n5098);
not gate_5072(n5100,n5099);
and gate_5073(n5101,n787,n5100);
not gate_5074(n5102,n5101);
and gate_5075(n5103,pi7,n5102);
not gate_5076(n5104,n5103);
and gate_5077(n5105,n45,n206);
not gate_5078(n5106,n5105);
and gate_5079(n5107,n5104,n5106);
not gate_5080(n5108,n5107);
and gate_5081(n5109,pi0,n5108);
not gate_5082(n5110,n5109);
and gate_5083(n5111,n45,n142);
not gate_5084(n5112,n5111);
and gate_5085(n5113,n5110,n5112);
and gate_5086(n5114,n5096,n5113);
not gate_5087(n5115,n5114);
and gate_5088(n5116,pi2,n5115);
not gate_5089(n5117,n5116);
and gate_5090(n5118,pi3,n181);
not gate_5091(n5119,n5118);
and gate_5092(n5120,n227,n4202);
not gate_5093(n5121,n5120);
and gate_5094(n5122,n5119,n5121);
not gate_5095(n5123,n5122);
and gate_5096(n5124,n2093,n5123);
not gate_5097(n5125,n5124);
and gate_5098(n5126,n5117,n5125);
not gate_5099(n5127,n5126);
and gate_5100(n5128,n31,n5127);
not gate_5101(n5129,n5128);
and gate_5102(n5130,n1234,n2571);
not gate_5103(n5131,n5130);
and gate_5104(n5132,n5129,n5131);
and gate_5105(n5133,n5082,n5132);
not gate_5106(n5134,n5133);
and gate_5107(n5135,pi5,n5134);
not gate_5108(n5136,n5135);
and gate_5109(n5137,n117,n163);
not gate_5110(n5138,n5137);
and gate_5111(n5139,pi1,n5138);
not gate_5112(n5140,n5139);
and gate_5113(n5141,n30,n5140);
not gate_5114(n5142,n5141);
and gate_5115(n5143,n801,n4488);
not gate_5116(n5144,n5143);
and gate_5117(n5145,n5142,n5144);
not gate_5118(n5146,n5145);
and gate_5119(n5147,n32,n5146);
not gate_5120(n5148,n5147);
and gate_5121(n5149,n5136,n5148);
and gate_5122(n5150,n5011,n5149);
not gate_5123(po14,n5150);
and gate_5124(n5152,n826,n1145);
not gate_5125(n5153,n5152);
and gate_5126(n5154,n299,n3116);
not gate_5127(n5155,n5154);
and gate_5128(n5156,n5153,n5155);
not gate_5129(n5157,n5156);
and gate_5130(n5158,pi4,n5157);
not gate_5131(n5159,n5158);
and gate_5132(n5160,n97,n299);
not gate_5133(n5161,n5160);
and gate_5134(n5162,n184,n1145);
not gate_5135(n5163,n5162);
and gate_5136(n5164,n5161,n5163);
not gate_5137(n5165,n5164);
and gate_5138(n5166,pi3,n5165);
not gate_5139(n5167,n5166);
and gate_5140(n5168,n51,n299);
not gate_5141(n5169,n5168);
and gate_5142(n5170,n5167,n5169);
not gate_5143(n5171,n5170);
and gate_5144(n5172,n34,n5171);
not gate_5145(n5173,n5172);
and gate_5146(n5174,n5159,n5173);
not gate_5147(n5175,n5174);
and gate_5148(n5176,pi5,n5175);
not gate_5149(n5177,n5176);
and gate_5150(n5178,n220,n2023);
and gate_5151(n5179,n299,n5178);
not gate_5152(n5180,n5179);
and gate_5153(n5181,n5177,n5180);
and gate_5154(n5182,n2149,n4761);
not gate_5155(n5183,n5182);
and gate_5156(n5184,n38,n5183);
not gate_5157(n5185,n5184);
and gate_5158(n5186,n31,n387);
not gate_5159(n5187,n5186);
and gate_5160(n5188,n5185,n5187);
not gate_5161(n5189,n5188);
and gate_5162(n5190,n37,n5189);
not gate_5163(n5191,n5190);
and gate_5164(n5192,n299,n1387);
not gate_5165(n5193,n5192);
and gate_5166(n5194,n5191,n5193);
not gate_5167(n5195,n5194);
and gate_5168(n5196,n36,n5195);
not gate_5169(n5197,n5196);
and gate_5170(n5198,pi4,n1274);
not gate_5171(n5199,n5198);
and gate_5172(n5200,pi1,n1270);
not gate_5173(n5201,n5200);
and gate_5174(n5202,n5199,n5201);
and gate_5175(n5203,n51,n5202);
and gate_5176(n5204,pi2,n5203);
not gate_5177(n5205,n5204);
and gate_5178(n5206,n5197,n5205);
not gate_5179(n5207,n5206);
and gate_5180(n5208,n35,n5207);
not gate_5181(n5209,n5208);
and gate_5182(n5210,n114,n1475);
not gate_5183(n5211,n5210);
and gate_5184(n5212,n143,n5211);
not gate_5185(n5213,n5212);
and gate_5186(n5214,n36,n5213);
not gate_5187(n5215,n5214);
and gate_5188(n5216,pi2,n5215);
not gate_5189(n5217,n5216);
and gate_5190(n5218,n31,n5217);
not gate_5191(n5219,n5218);
and gate_5192(n5220,n2064,n4760);
not gate_5193(n5221,n5220);
and gate_5194(n5222,n5219,n5221);
and gate_5195(n5223,n5209,n5222);
and gate_5196(n5224,n5181,n5223);
not gate_5197(n5225,n5224);
and gate_5198(po15,n30,n5225);
and gate_5199(n5227,n642,n1642);
not gate_5200(n5228,n5227);
and gate_5201(n5229,n31,n1192);
and gate_5202(n5230,n644,n5229);
not gate_5203(n5231,n5230);
and gate_5204(n5232,n5228,n5231);
and gate_5205(n5233,n181,n277);
and gate_5206(n5234,n4760,n5233);
not gate_5207(n5235,n5234);
and gate_5208(n5236,pi6,n583);
not gate_5209(n5237,n5236);
and gate_5210(n5238,n1752,n5237);
not gate_5211(n5239,n5238);
and gate_5212(n5240,n1166,n5239);
not gate_5213(n5241,n5240);
and gate_5214(n5242,n5235,n5241);
and gate_5215(n5243,n5232,n5242);
not gate_5216(n5244,n5243);
and gate_5217(n5245,n38,n5244);
not gate_5218(n5246,n5245);
and gate_5219(n5247,pi1,n1187);
not gate_5220(n5248,n5247);
and gate_5221(n5249,n4966,n5248);
not gate_5222(n5250,n5249);
and gate_5223(n5251,n35,n5250);
not gate_5224(n5252,n5251);
and gate_5225(n5253,n299,n509);
not gate_5226(n5254,n5253);
and gate_5227(n5255,n5252,n5254);
not gate_5228(n5256,n5255);
and gate_5229(n5257,n37,n5256);
not gate_5230(n5258,n5257);
and gate_5231(n5259,n1455,n5258);
not gate_5232(n5260,n5259);
and gate_5233(n5261,pi8,n5260);
not gate_5234(n5262,n5261);
and gate_5235(n5263,n299,n608);
not gate_5236(n5264,n5263);
and gate_5237(n5265,n5262,n5264);
not gate_5238(n5266,n5265);
and gate_5239(n5267,pi6,n5266);
not gate_5240(n5268,n5267);
and gate_5241(n5269,pi2,n257);
not gate_5242(n5270,n5269);
and gate_5243(n5271,n82,n5270);
not gate_5244(n5272,n5271);
and gate_5245(n5273,n35,n5272);
not gate_5246(n5274,n5273);
and gate_5247(n5275,pi4,n5274);
not gate_5248(n5276,n5275);
and gate_5249(n5277,n1155,n5276);
not gate_5250(n5278,n5277);
and gate_5251(n5279,n5268,n5278);
not gate_5252(n5280,n5279);
and gate_5253(n5281,n33,n5280);
not gate_5254(n5282,n5281);
and gate_5255(n5283,n1242,n5282);
and gate_5256(n5284,n5246,n5283);
not gate_5257(n5285,n5284);
and gate_5258(po16,n30,n5285);
and gate_5259(n5287,pi5,n5111);
not gate_5260(n5288,n5287);
and gate_5261(n5289,pi3,n155);
not gate_5262(n5290,n5289);
and gate_5263(n5291,n51,n1789);
not gate_5264(n5292,n5291);
and gate_5265(n5293,n5290,n5292);
not gate_5266(n5294,n5293);
and gate_5267(n5295,pi4,n5294);
not gate_5268(n5296,n5295);
and gate_5269(n5297,pi1,n5296);
and gate_5270(n5298,n5288,n5297);
not gate_5271(n5299,n5298);
and gate_5272(n5300,n32,n5299);
not gate_5273(n5301,n5300);
and gate_5274(n5302,n617,n2100);
not gate_5275(n5303,n5302);
and gate_5276(n5304,n257,n2162);
not gate_5277(n5305,n5304);
and gate_5278(n5306,n34,n695);
not gate_5279(n5307,n5306);
and gate_5280(n5308,n5305,n5307);
not gate_5281(n5309,n5308);
and gate_5282(n5310,n51,n5309);
not gate_5283(n5311,n5310);
and gate_5284(n5312,n5303,n5311);
not gate_5285(n5313,n5312);
and gate_5286(n5314,pi2,n5313);
not gate_5287(n5315,n5314);
and gate_5288(n5316,n787,n5315);
not gate_5289(n5317,n5316);
and gate_5290(n5318,n31,n5317);
not gate_5291(n5319,n5318);
and gate_5292(n5320,n5301,n5319);
not gate_5293(n5321,n5320);
and gate_5294(po17,n30,n5321);
and gate_5295(n5323,n104,n2870);
not gate_5296(n5324,n5323);
and gate_5297(n5325,n1325,n5324);
not gate_5298(n5326,n5325);
and gate_5299(n5327,n33,n5326);
not gate_5300(n5328,n5327);
and gate_5301(n5329,n627,n645);
not gate_5302(n5330,n5329);
and gate_5303(n5331,n1192,n5330);
not gate_5304(n5332,n5331);
and gate_5305(n5333,n5328,n5332);
not gate_5306(n5334,n5333);
and gate_5307(n5335,n35,n5334);
not gate_5308(n5336,n5335);
and gate_5309(n5337,n1954,n2908);
and gate_5310(n5338,pi2,n5337);
not gate_5311(n5339,n5338);
and gate_5312(n5340,n5336,n5339);
not gate_5313(n5341,n5340);
and gate_5314(n5342,n31,n5341);
not gate_5315(n5343,n5342);
and gate_5316(n5344,pi3,n3852);
not gate_5317(n5345,n5344);
and gate_5318(n5346,n3854,n5345);
and gate_5319(n5347,pi6,n5346);
not gate_5320(n5348,n5347);
and gate_5321(n5349,n258,n1006);
and gate_5322(n5350,n309,n5349);
not gate_5323(n5351,n5350);
and gate_5324(n5352,n5348,n5351);
not gate_5325(n5353,n5352);
and gate_5326(n5354,n1145,n5353);
not gate_5327(n5355,n5354);
and gate_5328(n5356,n5343,n5355);
not gate_5329(n5357,n5356);
and gate_5330(n5358,n38,n5357);
not gate_5331(n5359,n5358);
and gate_5332(n5360,n918,n1490);
and gate_5333(n5361,n1145,n5360);
not gate_5334(n5362,n5361);
and gate_5335(n5363,n88,n1168);
not gate_5336(n5364,n5363);
and gate_5337(n5365,n4965,n5364);
not gate_5338(n5366,n5365);
and gate_5339(n5367,n5362,n5366);
not gate_5340(n5368,n5367);
and gate_5341(n5369,pi8,n5368);
not gate_5342(n5370,n5369);
and gate_5343(n5371,pi1,n907);
and gate_5344(n5372,n996,n5371);
not gate_5345(n5373,n5372);
and gate_5346(n5374,n5370,n5373);
not gate_5347(n5375,n5374);
and gate_5348(n5376,pi3,n5375);
not gate_5349(n5377,n5376);
and gate_5350(n5378,n142,n146);
not gate_5351(n5379,n5378);
and gate_5352(n5380,pi2,n5379);
not gate_5353(n5381,n5380);
and gate_5354(n5382,n31,n5381);
not gate_5355(n5383,n5382);
and gate_5356(n5384,n5377,n5383);
and gate_5357(n5385,n5359,n5384);
not gate_5358(n5386,n5385);
and gate_5359(po18,n30,n5386);
endmodule
