// Verilog File 
module c7552 (G1,G5,G9,G12,G15,G18,G23,G26,G29,
G32,G35,G38,G41,G44,G47,G50,G53,G54,G55,
G56,G57,G58,G59,G60,G61,G62,G63,G64,G65,
G66,G69,G70,G73,G74,G75,G76,G77,G78,G79,
G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,
G94,G97,G100,G103,G106,G109,G110,G111,G112,G113,
G114,G115,G118,G121,G124,G127,G130,G133,G134,G135,
G138,G141,G144,G147,G150,G151,G152,G153,G154,G155,
G156,G157,G158,G159,G160,G161,G162,G163,G164,G165,
G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,
G176,G177,G178,G179,G180,G181,G182,G183,G184,G185,
G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,
G196,G197,G198,G199,G200,G201,G202,G203,G204,G205,
G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,
G216,G217,G218,G219,G220,G221,G222,G223,G224,G225,
G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,
G236,G237,G238,G239,G240,G1197,G1455,G1459,G1462,G1469,
G1480,G1486,G1492,G1496,G2204,G2208,G2211,G2218,G2224,G2230,
G2236,G2239,G2247,G2253,G2256,G3698,G3701,G3705,G3711,G3717,
G3723,G3729,G3737,G3743,G3749,G4393,G4394,G4400,G4405,G4410,
G4415,G4420,G4427,G4432,G4437,G4526,G4528,G2,G3,G450,
G448,G444,G442,G440,G438,G496,G494,G492,G490,G488,
G486,G484,G482,G480,G560,G542,G558,G556,G554,G552,
G550,G548,G546,G544,G540,G538,G536,G534,G532,G530,
G528,G526,G524,G279,G436,G478,G522,G402,G404,G406,
G408,G410,G432,G446,G284,G286,G289,G292,G341,G281,
G453,G278,G373,G246,G258,G264,G270,G388,G391,G394,
G397,G376,G379,G382,G385,G412,G414,G416,G249,G295,
G324,G252,G276,G310,G313,G316,G319,G327,G330,G333,
G336,G418,G273,G298,G301,G304,G307,G344,G422,G469,
G419,G471,G359,G362,G365,G368,G347,G350,G353,G356,
G321,G338,G370,G399);

input G1,G5,G9,G12,G15,G18,G23,G26,G29,
G32,G35,G38,G41,G44,G47,G50,G53,G54,G55,
G56,G57,G58,G59,G60,G61,G62,G63,G64,G65,
G66,G69,G70,G73,G74,G75,G76,G77,G78,G79,
G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,
G94,G97,G100,G103,G106,G109,G110,G111,G112,G113,
G114,G115,G118,G121,G124,G127,G130,G133,G134,G135,
G138,G141,G144,G147,G150,G151,G152,G153,G154,G155,
G156,G157,G158,G159,G160,G161,G162,G163,G164,G165,
G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,
G176,G177,G178,G179,G180,G181,G182,G183,G184,G185,
G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,
G196,G197,G198,G199,G200,G201,G202,G203,G204,G205,
G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,
G216,G217,G218,G219,G220,G221,G222,G223,G224,G225,
G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,
G236,G237,G238,G239,G240,G1197,G1455,G1459,G1462,G1469,
G1480,G1486,G1492,G1496,G2204,G2208,G2211,G2218,G2224,G2230,
G2236,G2239,G2247,G2253,G2256,G3698,G3701,G3705,G3711,G3717,
G3723,G3729,G3737,G3743,G3749,G4393,G4394,G4400,G4405,G4410,
G4415,G4420,G4427,G4432,G4437,G4526,G4528;

output G2,G3,G450,G448,G444,G442,G440,G438,G496,
G494,G492,G490,G488,G486,G484,G482,G480,G560,G542,
G558,G556,G554,G552,G550,G548,G546,G544,G540,G538,
G536,G534,G532,G530,G528,G526,G524,G279,G436,G478,
G522,G402,G404,G406,G408,G410,G432,G446,G284,G286,
G289,G292,G341,G281,G453,G278,G373,G246,G258,G264,
G270,G388,G391,G394,G397,G376,G379,G382,G385,G412,
G414,G416,G249,G295,G324,G252,G276,G310,G313,G316,
G319,G327,G330,G333,G336,G418,G273,G298,G301,G304,
G307,G344,G422,G469,G419,G471,G359,G362,G365,G368,
G347,G350,G353,G356,G321,G338,G370,G399;

wire G400,G1184,G1501,G2857,G4442,G4514,G401,G573,G574,
G575,G1178,G1186,G1192,G1198,G1205,G1206,G1207,G1210,G1458,
G1461,G1464,G1471,G1475,G1482,G1488,G1495,G1499,G1500,G1503,
G1512,G1518,G1524,G1535,G1541,G2207,G2210,G2213,G2220,G2226,
G2232,G2238,G2241,G2249,G2255,G2258,G2828,G3700,G3703,G3707,
G3713,G3719,G3725,G3731,G3739,G3745,G3751,G4121,G4396,G4402,
G4407,G4412,G4417,G4422,G4429,G4434,G4439,G4833,G2876,G2878,
G1519,G2871,G2883,G280,G4839,G572,G581,G587,G601,G606,
G650,G657,G671,G678,G777,G1115,G1336,G1350,G1477,G1507,
G1514,G1530,G2259,G2833,G2872,G2886,G2892,G2905,G2909,G3622,
G3635,G3755,G4640,G4653,G4873,G4876,G4881,G4889,G4905,G4916,
G4921,G5175,G5178,G5186,G5191,G5199,G5215,G5223,G5393,G5401,
G5409,G5417,G5425,G5433,G5441,G5449,G5457,G5745,G5753,G5761,
G5769,G5777,G5785,G5793,G5801,G5809,G5865,G5873,G5881,G5889,
G5897,G5905,G5913,G5921,G5985,G5993,G6001,G6009,G6017,G6025,
G6033,G6041,G6514,G6554,G6567,G6575,G6583,G6591,G6599,G6607,
G6615,G6623,G6631,G6853,G6861,G6869,G6877,G6885,G6893,G6901,
G6909,G6917,G784,G1014,G3221,G4913,G4929,G5183,G5231,G6511,
G615,G594,G611,G617,G619,G621,G623,G625,G627,G664,
G685,G691,G693,G695,G697,G699,G701,G703,G705,G707,
G709,G4879,G4880,G4887,G4895,G4911,G4920,G4927,G5181,G5182,
G5190,G5197,G5205,G5221,G5229,G1343,G1357,G1364,G1366,G1368,
G1370,G1372,G1374,G1376,G1378,G1380,G1382,G5399,G5407,G5415,
G5423,G5431,G5439,G5447,G5455,G5463,G5751,G5759,G5767,G5775,
G5783,G5791,G5799,G5807,G5815,G2019,G2032,G2117,G2130,G2266,
G2272,G2286,G2288,G2290,G2292,G2294,G5871,G5879,G5887,G5895,
G5903,G5911,G5919,G5927,G5991,G5999,G6007,G6015,G6023,G6031,
G6039,G6047,G2899,G2914,G2919,G2921,G2923,G2925,G2927,G2929,
G2931,G6518,G3173,G6558,G6573,G6581,G6589,G6597,G6605,G6613,
G6621,G6629,G6637,G3629,G3642,G3649,G3651,G3653,G3655,G3657,
G3659,G3661,G3663,G3762,G3768,G3782,G3784,G3786,G3788,G3790,
G6859,G6867,G6875,G6883,G6891,G6899,G6907,G6915,G6923,G4094,
G4107,G4444,G4457,G4647,G4660,G4667,G4669,G4671,G4673,G4675,
G4677,G4679,G4681,G4683,G4685,G4897,G5207,G6551,G763,G764,
G4919,G886,G1005,G1006,G5189,G1018,G5237,G6517,G3169,G4935,
G4970,G5239,G577,G616,G618,G620,G622,G624,G626,G628,
G692,G694,G696,G698,G700,G702,G704,G706,G708,G710,
G765,G4903,G885,G1007,G1017,G5213,G1363,G1365,G1367,G1369,
G1371,G1373,G1375,G1377,G1379,G1381,G2026,G2039,G2046,G2048,
G2050,G2052,G2054,G2056,G2058,G2060,G2062,G2064,G2124,G2137,
G2144,G2146,G2148,G2150,G2152,G2154,G2156,G2158,G2160,G2162,
G2279,G2285,G2287,G2289,G2291,G2293,G2296,G2298,G2300,G2302,
G2304,G2918,G2920,G2922,G2924,G2926,G2928,G2930,G2932,G3168,
G6557,G3211,G3648,G3650,G3652,G3654,G3656,G3658,G3660,G3662,
G3665,G3666,G3775,G3781,G3783,G3785,G3787,G3789,G3792,G3794,
G3796,G3798,G3800,G4101,G4114,G4123,G4126,G4129,G4132,G4135,
G4138,G4141,G4144,G4147,G4150,G4451,G4464,G4471,G4473,G4475,
G4477,G4479,G4481,G4483,G4485,G4487,G4489,G4666,G4668,G4670,
G4672,G4674,G4676,G4678,G4680,G4682,G4684,G579,G629,G633,
G637,G641,G645,G711,G715,G719,G723,G727,G731,G737,
G745,G751,G757,G887,G1019,G5245,G1383,G1387,G1391,G1395,
G1399,G1406,G1412,G1418,G2305,G2308,G2312,G2316,G2933,G2938,
G2942,G2946,G2950,G3170,G3210,G3667,G3670,G3673,G3676,G3679,
G3682,G3686,G3801,G3804,G3807,G3810,G3813,G4525,G4686,G4689,
G4692,G4695,G4698,G4701,G4704,G4707,G4710,G4976,G5271,G5274,
G5305,G5308,G5318,G6690,G6711,G6714,G7252,G7296,G7466,G907,
G913,G915,G916,G1116,G2045,G2047,G2049,G2051,G2053,G2055,
G2057,G2059,G2061,G2063,G2143,G2145,G2147,G2149,G2151,G2153,
G2155,G2157,G2159,G2161,G2295,G2297,G2299,G2301,G2303,G3212,
G3791,G3793,G3795,G3797,G3799,G4122,G4125,G4128,G4131,G4134,
G4137,G4140,G4143,G4146,G4149,G4470,G4472,G4474,G4476,G4478,
G4480,G4482,G4484,G4486,G4488,G4962,G5003,G5234,G5242,G5250,
G5284,G802,G821,G845,G868,G877,G902,G908,G914,G917,
G953,G1023,G1035,G1050,G1068,G1086,G1102,G1108,G1117,G5322,
G1553,G1567,G1584,G1590,G1606,G1624,G1647,G1669,G1677,G1802,
G1816,G1834,G1841,G1866,G1880,G1897,G1914,G1929,G2065,G2069,
G2073,G2077,G2081,G2085,G2091,G2099,G2105,G2111,G2163,G2167,
G2171,G2175,G2179,G2186,G2192,G2198,G2320,G2323,G2329,G2335,
G2962,G2970,G2977,G2979,G2989,G2998,G3006,G3013,G3015,G3183,
G3192,G3200,G3207,G3209,G3216,G3222,G6694,G3695,G3816,G3821,
G3828,G3833,G3838,G4151,G4154,G4157,G4160,G4163,G4166,G4169,
G4172,G4175,G7256,G7300,G4490,G4493,G4496,G4499,G4502,G4505,
G4508,G4511,G7470,G4884,G4892,G4900,G4908,G4924,G4952,G4983,
G4993,G5011,G5194,G5202,G5210,G5218,G5226,G5247,G5255,G5258,
G5263,G5266,G5277,G5278,G5281,G5289,G5292,G5297,G5300,G5311,
G5312,G5315,G5323,G5326,G5331,G5334,G5339,G5342,G5349,G5352,
G5396,G5404,G5412,G5420,G5428,G5436,G5444,G5452,G5460,G5465,
G5581,G5748,G5756,G5764,G5772,G5780,G5788,G5796,G5804,G5812,
G5849,G5929,G6049,G6367,G6370,G6375,G6378,G6383,G6386,G6391,
G6394,G6399,G6402,G6407,G6410,G6415,G6418,G6423,G6426,G6431,
G6434,G6442,G6450,G6458,G6466,G6498,G6519,G6522,G6527,G6530,
G6535,G6538,G6543,G6546,G6559,G6562,G6687,G6695,G6698,G6703,
G6706,G6717,G6718,G6724,G6768,G7208,G7221,G7229,G7232,G7239,
G7242,G7249,G7257,G7260,G7268,G7293,G7301,G7304,G7309,G7312,
G7317,G7320,G7327,G7330,G7396,G7404,G7412,G7425,G7463,G7471,
G7474,G7479,G7482,G7487,G7490,G7497,G7500,G7507,G7510,G7554,
G1152,G5238,G1156,G5246,G5254,G5288,G3223,G4942,G4966,G5007,
G5279,G5280,G5313,G5314,G6719,G6720,G790,G4888,G803,G4896,
G825,G4904,G851,G4912,G893,G4928,G906,G912,G1024,G5198,
G1036,G5206,G1053,G5214,G1072,G5222,G1091,G5230,G1112,G1121,
G1153,G1157,G5253,G1216,G5261,G5262,G5269,G5270,G5287,G1239,
G5295,G5296,G5303,G5304,G5321,G1262,G5329,G5330,G5337,G5338,
G1544,G5400,G1554,G5408,G1571,G5416,G1596,G5424,G1607,G5432,
G1628,G5440,G1653,G5448,G1685,G5456,G1693,G5464,G1793,G5752,
G1803,G5760,G1820,G5768,G1848,G5776,G1857,G5784,G1867,G5792,
G1883,G5800,G1901,G5808,G1919,G5816,G5855,G2351,G2366,G2384,
G2391,G2417,G2431,G2448,G2465,G5935,G2597,G2612,G2629,G2635,
G2652,G2670,G2693,G2715,G6055,G6373,G6374,G6381,G6382,G6389,
G6390,G6397,G6398,G6405,G6406,G6413,G6414,G6421,G6422,G6429,
G6430,G6437,G6438,G6446,G3059,G6454,G3068,G6462,G3076,G3079,
G6470,G3090,G3099,G3107,G3114,G3116,G6502,G6525,G6526,G6533,
G6534,G6541,G6542,G6549,G6550,G6565,G6566,G3220,G3292,G3308,
G3327,G3335,G3362,G3376,G3393,G3410,G3425,G6693,G3503,G6701,
G6702,G6709,G6710,G6728,G6772,G3853,G3868,G3885,G3891,G3908,
G3926,G3949,G3971,G3979,G7212,G7227,G7255,G4202,G7263,G7264,
G7272,G7299,G4225,G7307,G7308,G7315,G7316,G4297,G4305,G4312,
G4314,G4324,G7400,G4333,G7408,G4341,G7416,G4348,G4349,G7431,
G4389,G7469,G4530,G7477,G7478,G7485,G7486,G7513,G7514,G7558,
G4932,G4956,G4973,G4987,G4997,G5017,G5099,G5345,G5346,G5355,
G5356,G5372,G5380,G5471,G5523,G5587,G5669,G5857,G5868,G5876,
G5884,G5892,G5900,G5908,G5916,G5924,G5969,G5988,G5996,G6004,
G6012,G6020,G6028,G6036,G6044,G6057,G6439,G6447,G6455,G6463,
G6471,G6474,G6479,G6482,G6487,G6490,G6495,G6503,G6506,G6570,
G6578,G6586,G6594,G6602,G6610,G6618,G6626,G6634,G6671,G6721,
G6729,G6732,G6737,G6740,G6745,G6748,G6755,G6758,G6765,G6773,
G6776,G6781,G6784,G6789,G6792,G6799,G6802,G6832,G6856,G6864,
G6872,G6880,G6888,G6896,G6904,G6912,G6920,G6925,G7041,G7205,
G7213,G7216,G7224,G7235,G7236,G7245,G7246,G7265,G7273,G7276,
G7283,G7286,G7323,G7324,G7333,G7334,G7361,G7364,G7369,G7372,
G7377,G7380,G7385,G7388,G7393,G7401,G7409,G7417,G7420,G7428,
G7493,G7494,G7503,G7504,G7515,G7518,G7523,G7526,G7531,G7534,
G7541,G7544,G7551,G7559,G7562,G7567,G7570,G7575,G7578,G7585,
G7588,G1176,G957,G791,G804,G826,G852,G894,G1025,G1037,
G1054,G1073,G1092,G1154,G1158,G1215,G1224,G1225,G1233,G1234,
G1238,G1247,G1248,G1256,G1257,G1261,G1270,G1271,G1279,G1280,
G1545,G1555,G1572,G1597,G1608,G1629,G1654,G1686,G1694,G1794,
G1804,G1821,G1849,G1858,G1868,G1884,G1902,G1920,G2954,G2955,
G2963,G2964,G2971,G2972,G2980,G2981,G2990,G2991,G2999,G3000,
G3007,G3008,G3016,G3017,G3019,G3020,G3174,G3175,G3184,G3185,
G3193,G3194,G3201,G3202,G3213,G3214,G3227,G3502,G3511,G3512,
G3520,G3521,G4201,G4210,G4211,G4224,G4233,G4234,G4242,G4243,
G4529,G4538,G4539,G4547,G4548,G4552,G4553,G4946,G5347,G5348,
G5357,G5358,G7237,G7238,G7247,G7248,G7325,G7326,G7335,G7336,
G7495,G7496,G7505,G7506,G3244,G792,G805,G827,G853,G895,
G1026,G1038,G1055,G1074,G1093,G1155,G1217,G1226,G1235,G1240,
G1249,G1258,G1263,G1272,G1281,G5376,G5384,G1546,G1556,G1573,
G1598,G1609,G1630,G1655,G1687,G1695,G1795,G1805,G1822,G1850,
G1859,G1869,G1885,G1903,G1921,G5863,G2341,G5872,G2352,G5880,
G2370,G5888,G2398,G5896,G2407,G5904,G2418,G5912,G2434,G5920,
G2452,G5928,G2481,G5975,G2587,G5992,G2598,G6000,G2616,G6008,
G2641,G6016,G2653,G6024,G2674,G6032,G2699,G6040,G2724,G2732,
G6048,G2956,G2965,G2973,G2982,G2992,G3001,G3009,G3018,G3021,
G6445,G3051,G6453,G3061,G6461,G3070,G6469,G3081,G6477,G6478,
G6485,G6486,G6493,G6494,G6501,G3118,G6509,G6510,G3176,G3186,
G3195,G3203,G3215,G3281,G6574,G3293,G6582,G3312,G6590,G3342,
G6598,G3351,G6606,G3363,G6614,G3379,G6622,G3397,G6630,G3415,
G6638,G6677,G3504,G3513,G3522,G6727,G3526,G6735,G6736,G6743,
G6744,G6771,G3549,G6779,G6780,G6787,G6788,G6836,G3843,G6860,
G3854,G6868,G3872,G6876,G3897,G6884,G3909,G6892,G3930,G6900,
G3955,G6908,G3987,G6916,G3995,G6924,G7211,G4179,G7219,G7220,
G4196,G7228,G4203,G4212,G7271,G4220,G4226,G4235,G4244,G7367,
G7368,G7375,G7376,G7383,G7384,G7391,G7392,G7399,G4326,G7407,
G4335,G7415,G4343,G7423,G7424,G4353,G7432,G4531,G4540,G4549,
G4554,G7521,G7522,G7529,G7530,G7557,G4576,G7565,G7566,G7573,
G7574,G4936,G4937,G4977,G4978,G5105,G5359,G5362,G5529,G5675,
G5932,G5977,G6052,G6063,G6115,G6173,G6679,G6751,G6752,G6761,
G6762,G6795,G6796,G6805,G6806,G6931,G6983,G7047,G7129,G7279,
G7280,G7289,G7290,G7337,G7340,G7353,G7356,G7537,G7538,G7547,
G7548,G7581,G7582,G7591,G7592,G7595,G7598,G2342,G2353,G2371,
G2399,G2408,G2419,G2435,G2453,G2588,G2599,G2617,G2642,G2654,
G2675,G2700,G2733,G3050,G3060,G3069,G3080,G3091,G3092,G3100,
G3101,G3108,G3109,G3117,G3120,G3121,G3282,G3294,G3313,G3343,
G3352,G3364,G3380,G3398,G3416,G3525,G3534,G3535,G3543,G3544,
G3548,G3557,G3558,G3566,G3567,G3844,G3855,G3873,G3898,G3910,
G3931,G3956,G3988,G3996,G4178,G4187,G4188,G4197,G4219,G4289,
G4290,G4298,G4299,G4306,G4307,G4315,G4316,G4325,G4334,G4342,
G4350,G4351,G4354,G4561,G4562,G4570,G4571,G4575,G4584,G4585,
G4593,G4594,G4938,G4979,G6753,G6754,G6763,G6764,G6797,G6798,
G6807,G6808,G7281,G7282,G7291,G7292,G7539,G7540,G7549,G7550,
G7583,G7584,G7593,G7594,G1856,G920,G925,G926,G927,G928,
G937,G938,G939,G940,G941,G942,G943,G944,G945,G946,
G947,G948,G949,G956,G1122,G1125,G1126,G1127,G1128,G1132,
G1133,G1134,G1137,G1138,G1141,G1221,G1230,G1244,G1253,G1267,
G1276,G1284,G1288,G1292,G1296,G1300,G1304,G1702,G1705,G1706,
G1707,G1709,G1710,G1711,G1712,G1713,G1714,G1718,G1722,G1723,
G1724,G1725,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1740,
G1741,G1742,G1743,G1744,G1745,G1749,G1750,G1935,G1938,G1939,
G1940,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,
G1953,G1954,G1955,G1956,G1960,G1961,G1962,G1965,G1966,G1969,
G2343,G2354,G2372,G2400,G2409,G2420,G2436,G2454,G2470,G5936,
G5983,G2589,G2600,G2618,G2643,G2655,G2676,G2701,G2734,G2740,
G6056,G3022,G3025,G3026,G3027,G3029,G3030,G3031,G3032,G3033,
G3052,G3062,G3071,G3082,G3093,G3102,G3110,G3119,G3122,G3228,
G3231,G3232,G3233,G3234,G3283,G3295,G3314,G3344,G3353,G3365,
G3381,G3399,G3417,G6685,G3508,G3517,G3527,G3536,G3545,G3550,
G3559,G3568,G3571,G3575,G3845,G3856,G3874,G3899,G3911,G3932,
G3957,G3989,G3997,G4180,G4189,G4198,G4207,G4216,G4221,G4230,
G4239,G4263,G4267,G4291,G4300,G4308,G4317,G4327,G4336,G4344,
G4352,G4355,G4535,G4544,G4558,G4563,G4572,G4577,G4586,G4595,
G4598,G4602,G4716,G4724,G4732,G4740,G4748,G4756,G4764,G4772,
G4780,G4788,G4939,G4980,G5044,G5054,G5064,G5074,G5084,G5094,
G5132,G5142,G5152,G5162,G5365,G5366,G5488,G5498,G5508,G5518,
G5546,G5556,G5566,G5576,G5614,G5624,G5634,G5644,G5654,G5664,
G5702,G5712,G5722,G5732,G5820,G5828,G5836,G5844,G5852,G5860,
G6121,G6179,G6261,G7359,G7360,G7343,G7344,G6809,G6812,G6819,
G6822,G6989,G7135,G7345,G7348,G7601,G7602,G7603,G7606,G7611,
G7614,G929,G950,G1129,G1708,G1715,G1726,G1746,G1941,G1957,
G2471,G2741,G3028,G3034,G3235,G5014,G5034,G5102,G5122,G5367,
G5368,G5478,G5536,G5584,G5604,G5672,G5692,G5817,G5825,G5833,
G5841,G6340,G6341,G6350,G6351,G7436,G7437,G4720,G4728,G4736,
G4744,G4752,G4760,G4768,G4776,G4784,G4792,G3350,G2406,G924,
G5088,G5098,G997,G1146,G1287,G1291,G1295,G1299,G1303,G1307,
G1309,G1312,G1315,G1318,G1321,G1324,G1721,G5522,G5580,G5658,
G5668,G1788,G1974,G5824,G5832,G5840,G5848,G1999,G5856,G2003,
G5864,G2472,G2487,G2492,G2493,G2494,G2500,G2501,G2502,G2503,
G2504,G2505,G2506,G2507,G2511,G2512,G2513,G2514,G2518,G2519,
G2520,G2523,G2524,G2527,G2742,G2749,G2754,G2755,G2756,G2762,
G2763,G2764,G2765,G2766,G2767,G2776,G2777,G2778,G2779,G2788,
G2789,G2790,G2792,G2793,G2794,G2795,G2796,G2798,G2799,G2800,
G2804,G3035,G3045,G3123,G3128,G3129,G3130,G3136,G3139,G3140,
G3141,G3142,G3249,G3431,G3434,G3435,G3436,G3438,G3439,G3440,
G3441,G3442,G3443,G3444,G3445,G3446,G3449,G3450,G3451,G3452,
G3456,G3457,G3458,G3460,G3461,G3463,G3531,G3540,G3554,G3563,
G3574,G3578,G3579,G3583,G3587,G3591,G3596,G3599,G4004,G4007,
G4008,G4009,G4011,G4012,G4013,G4014,G4015,G4016,G4020,G4024,
G4025,G4026,G4027,G4035,G4036,G4037,G4038,G4039,G4040,G4041,
G4042,G4043,G4044,G4045,G4046,G4047,G4051,G4052,G4184,G4193,
G4247,G4251,G4255,G4259,G4266,G4270,G4284,G4287,G4356,G4361,
G4362,G4363,G4369,G4372,G4373,G4374,G4375,G4567,G4581,G4590,
G4601,G4605,G4606,G4610,G4614,G4618,G4623,G4626,G4796,G4804,
G4812,G4820,G4828,G4844,G4852,G4860,G4868,G4945,G4948,G4986,
G4989,G5048,G5058,G5068,G5078,G5166,G5136,G5146,G5156,G5388,
G5492,G5502,G5512,G5550,G5560,G5570,G5618,G5628,G5638,G5648,
G5736,G5706,G5716,G5726,G5940,G5948,G5956,G5964,G5972,G5980,
G6080,G6090,G6100,G6110,G6138,G6148,G6158,G6168,G6216,G6226,
G6236,G6246,G6256,G6267,G6304,G6314,G6324,G6342,G6352,G7351,
G7352,G6642,G6650,G6658,G6666,G6674,G6682,G6815,G6816,G6825,
G6826,G6948,G6958,G6968,G6978,G7006,G7016,G7026,G7036,G7074,
G7084,G7094,G7104,G7114,G7124,G7162,G7172,G7182,G7192,G7438,
G7617,G7618,G7609,G7610,G1151,G1002,G933,G1308,G1311,G1314,
G1317,G1320,G1323,G1730,G1789,G1981,G5823,G1986,G5831,G1989,
G5839,G1993,G5847,G1996,G2000,G2004,G2495,G2515,G2757,G2768,
G2780,G2801,G3046,G3131,G3143,G3238,G3258,G3437,G3453,G3595,
G3598,G4010,G4017,G4028,G4048,G4283,G4286,G4364,G4376,G4622,
G4625,G4947,G4988,G5018,G5019,G5024,G5038,G5106,G5107,G5112,
G5126,G5468,G5482,G5526,G5540,G5588,G5589,G5594,G5608,G5676,
G5677,G5682,G5696,G5937,G5945,G5953,G5961,G6070,G6128,G6264,
G6284,G6360,G6361,G6639,G6647,G6655,G6663,G6817,G6818,G6827,
G6828,G6938,G6996,G7044,G7064,G7132,G7152,G7446,G7447,G7456,
G7457,G241,G265,G2005,G4800,G4808,G4816,G4824,G4832,G4848,
G4856,G4864,G4872,G1310,G1313,G1316,G1319,G1322,G1325,G5392,
G1790,G1982,G1985,G1988,G1992,G1995,G2001,G2491,G2508,G2522,
G2526,G2529,G2531,G5944,G5952,G5960,G5968,G2555,G5976,G2559,
G5984,G2753,G2771,G2791,G2797,G2807,G6114,G6172,G6250,G6260,
G6346,G6356,G3127,G3156,G3259,G3466,G6646,G6654,G6662,G6670,
G3483,G6678,G3487,G6686,G3582,G3586,G3590,G3594,G3597,G3600,
G3602,G3605,G3608,G3611,G4023,G6982,G7040,G7118,G7128,G4089,
G4250,G4254,G4258,G4262,G4272,G4275,G4278,G4281,G4285,G4288,
G4360,G4380,G4386,G7442,G4609,G4613,G4617,G4621,G4624,G4627,
G4629,G4632,G4635,G4638,G4836,G4949,G4990,G5020,G5108,G5590,
G5678,G6084,G6094,G6104,G6142,G6152,G6162,G6206,G6220,G6230,
G6240,G6328,G6294,G6308,G6318,G6362,G6840,G6848,G6952,G6962,
G6972,G7010,G7020,G7030,G7078,G7088,G7098,G7108,G7196,G7166,
G7176,G7186,G7448,G7458,G254,G260,G1987,G1994,G2002,G962,
G1751,G1990,G1997,G2499,G2536,G5943,G2542,G5951,G2545,G5959,
G2549,G5967,G2552,G2556,G2560,G2761,G2784,G2853,G3135,G3146,
G3163,G3467,G6645,G3470,G6653,G3473,G6661,G3477,G6669,G3480,
G3484,G3488,G3601,G3604,G3607,G3610,G4032,G4090,G4271,G4274,
G4277,G4280,G4368,G4379,G4387,G4628,G4631,G4634,G4637,G4841,
G4849,G4857,G4865,G5021,G5028,G5109,G5116,G5369,G5377,G5385,
G5472,G5473,G5530,G5531,G5591,G5598,G5679,G5686,G6060,G6074,
G6118,G6132,G6176,G6186,G6196,G6268,G6269,G6274,G6288,G6337,
G6829,G6928,G6942,G6986,G7000,G7048,G7049,G7054,G7068,G7136,
G7137,G7142,G7156,G7433,G242,G3151,G257,G263,G266,G1991,
G1998,G3489,G371,G4840,G2561,G2532,G2537,G2541,G2544,G2548,
G2551,G2557,G2563,G2577,G2775,G2806,G2808,G2852,G2854,G6366,
G4381,G3164,G3241,G3468,G3469,G3472,G3476,G3479,G3485,G3603,
G3606,G3609,G3612,G6844,G6852,G4091,G4273,G4276,G4279,G4282,
G4382,G4388,G7452,G7462,G4630,G4633,G4636,G4639,G4955,G4958,
G4996,G4999,G5474,G5532,G6210,G6270,G6298,G7050,G7138,G3471,
G3478,G3486,G372,G2543,G2550,G2558,G4847,G387,G4855,G390,
G4863,G393,G4871,G396,G965,G5375,G1327,G5383,G1330,G5391,
G1333,G1754,G2546,G2553,G2564,G2809,G2813,G6345,G2860,G3474,
G3481,G6835,G3614,G4053,G7441,G4516,G4957,G4998,G5027,G5030,
G5115,G5118,G5475,G5533,G5597,G5600,G5685,G5688,G6064,G6065,
G6122,G6123,G6180,G6181,G6190,G6200,G6271,G6278,G6347,G6357,
G6837,G6845,G6932,G6933,G6990,G6991,G7051,G7058,G7139,G7146,
G7443,G7453,G243,G244,G245,G255,G256,G261,G262,G267,
G268,G269,G3475,G3482,G2547,G2554,G386,G389,G392,G395,
G1326,G1329,G1332,G1436,G1440,G1445,G1450,G1454,G2859,G4385,
G3148,G3239,G3240,G3265,G3267,G3270,G3274,G3277,G3613,G4515,
G4959,G5000,G5029,G5117,G5599,G5687,G6066,G6124,G6182,G6934,
G6992,G375,G378,G381,G384,G1328,G1331,G1334,G1447,G1766,
G2571,G2579,G2812,G2816,G2851,G2861,G6355,G2863,G6365,G2866,
G3147,G3242,G3271,G3279,G3615,G6843,G3617,G6851,G3620,G4056,
G4517,G7451,G4519,G7461,G4522,G5031,G5119,G5481,G5484,G5539,
G5542,G5601,G5689,G6067,G6125,G6183,G6277,G6280,G6935,G6993,
G7057,G7060,G7145,G7148,G4968,G5009,G2850,G2862,G2865,G3149,
G3243,G3616,G3619,G4518,G4521,G4965,G5006,G5483,G5541,G6279,
G7059,G7147,G374,G377,G380,G383,G955,G4967,G5008,G975,
G1136,G1140,G1143,G1145,G1160,G1771,G1964,G1968,G1971,G1973,
G2007,G2578,G2864,G2867,G3150,G3245,G3618,G3621,G4067,G4520,
G4523,G4713,G4753,G5037,G5040,G5125,G5128,G5485,G5543,G5607,
G5610,G5695,G5698,G6073,G6076,G6131,G6134,G6189,G6192,G6281,
G6941,G6944,G6999,G7002,G7061,G7149,G958,G967,G971,G1161,
G2008,G2580,G2868,G3152,G4443,G4524,G4721,G4729,G4737,G4745,
G4761,G4769,G4777,G4785,G5039,G5127,G5609,G5697,G6075,G6133,
G6191,G6943,G7001,G3248,G248,G4719,G294,G4759,G323,G980,
G4072,G5041,G5129,G5491,G5494,G5549,G5552,G5611,G5699,G6077,
G6135,G6193,G6287,G6290,G6945,G7003,G7067,G7070,G7155,G7158,
G247,G3155,G251,G272,G961,G275,G293,G297,G300,G303,
G306,G4727,G309,G4735,G312,G4743,G315,G4751,G318,G322,
G4767,G326,G4775,G329,G4783,G332,G4791,G335,G2881,G993,
G994,G1166,G1171,G1174,G2014,G3459,G3462,G3464,G3465,G3490,
G4793,G5493,G5551,G6289,G7069,G7157,G250,G274,G308,G311,
G314,G317,G325,G328,G331,G334,G417,G991,G992,G3491,
G4801,G4809,G4817,G4825,G5047,G5050,G5135,G5138,G5495,G5553,
G5617,G5620,G5705,G5708,G6083,G6086,G6141,G6144,G6199,G6202,
G6291,G6951,G6954,G7009,G7012,G7071,G7159,G271,G296,G299,
G302,G305,G4799,G343,G1170,G1173,G5049,G5137,G5167,G5619,
G5707,G6085,G6143,G6201,G6953,G7011,G342,G346,G349,G352,
G355,G4807,G358,G4815,G361,G4823,G364,G4831,G367,G1172,
G1175,G3497,G5051,G5139,G5501,G5504,G5559,G5562,G5621,G5709,
G6087,G6145,G6203,G6297,G6300,G6955,G7013,G7077,G7080,G7165,
G7168,G357,G360,G363,G366,G5173,G5503,G5561,G6299,G7079,
G7167,G345,G348,G351,G354,G5057,G5060,G5145,G5148,G5505,
G5563,G5627,G5630,G5715,G5718,G6093,G6096,G6151,G6154,G6209,
G6212,G6301,G6961,G6964,G7019,G7022,G7081,G7169,G5059,G5147,
G5629,G5717,G6095,G6153,G6211,G6963,G7021,G5061,G5149,G5511,
G5514,G5569,G5572,G5631,G5719,G6097,G6155,G6213,G6307,G6310,
G6965,G7023,G7087,G7090,G7175,G7178,G5513,G5571,G6309,G7089,
G7177,G5067,G5070,G5155,G5158,G5515,G5573,G5637,G5640,G5725,
G5728,G6103,G6106,G6161,G6164,G6219,G6222,G6311,G6971,G6974,
G7029,G7032,G7091,G7179,G5069,G5157,G5639,G5727,G6105,G6163,
G6221,G6973,G7031,G5521,G1756,G5579,G1761,G5071,G5159,G5641,
G5729,G6107,G6165,G6223,G6317,G6320,G6975,G7033,G7097,G7100,
G7185,G7188,G1755,G1760,G6319,G7099,G7187,G1757,G1762,G6113,
G2818,G6171,G2823,G6981,G4058,G7039,G4063,G5077,G5080,G5165,
G5090,G5647,G5650,G5735,G5660,G6229,G6232,G6321,G7101,G7189,
G2817,G2822,G4057,G4062,G5079,G5089,G5649,G5659,G6231,G1782,
G1783,G1784,G1785,G2819,G2824,G4059,G4064,G5081,G5091,G5651,
G5661,G6233,G6327,G6252,G7107,G7110,G7195,G7120,G5737,G6251,
G7109,G7119,G5087,G985,G5097,G988,G5657,G1776,G5667,G1779,
G2844,G2845,G2846,G2847,G4083,G4084,G4085,G4086,G6239,G6242,
G6253,G7111,G7121,G984,G987,G1775,G1778,G5743,G6241,G6329,
G7197,G986,G989,G1777,G1780,G6259,G2841,G7117,G4077,G7127,
G4080,G6243,G990,G996,G1781,G1787,G2840,G6335,G4076,G4079,
G7203,G995,G1786,G6249,G2838,G2842,G4078,G4081,G2837,G2843,
G4082,G4088,G5170,G5740,G2839,G2848,G4087,G1791,G1003,G5174,
G5744,G2849,G7200,G1792,G1004,G6332,G320,G337,G4092,G7204,
G4093,G2855,G6336,G369,G2856,G398;
buf gate_0(G2,G1);
buf gate_1(G3,G1);
not gate_2(G400,G57);
and gate_3(G1184,G134,G133);
buf gate_4(G450,G1459);
buf gate_5(G448,G1469);
buf gate_6(G444,G1480);
buf gate_7(G442,G1486);
buf gate_8(G440,G1492);
buf gate_9(G438,G1496);
and gate_10(G1501,G162,G172,G188,G199);
buf gate_11(G496,G2208);
buf gate_12(G494,G2218);
buf gate_13(G492,G2224);
buf gate_14(G490,G2230);
buf gate_15(G488,G2236);
buf gate_16(G486,G2239);
buf gate_17(G484,G2247);
buf gate_18(G482,G2253);
buf gate_19(G480,G2256);
and gate_20(G2857,G150,G184,G228,G240);
buf gate_21(G560,G3698);
buf gate_22(G542,G3701);
buf gate_23(G558,G3705);
buf gate_24(G556,G3711);
buf gate_25(G554,G3717);
buf gate_26(G552,G3723);
buf gate_27(G550,G3729);
buf gate_28(G548,G3737);
buf gate_29(G546,G3743);
buf gate_30(G544,G3749);
buf gate_31(G540,G4393);
buf gate_32(G538,G4400);
buf gate_33(G536,G4405);
buf gate_34(G534,G4410);
buf gate_35(G532,G4415);
buf gate_36(G530,G4420);
buf gate_37(G528,G4427);
buf gate_38(G526,G4432);
buf gate_39(G524,G4437);
and gate_40(G4442,G183,G182,G185,G186);
and gate_41(G4514,G210,G152,G218,G230);
not gate_42(G279,G15);
not gate_43(G401,G5);
buf gate_44(G573,G1);
not gate_45(G574,G5);
not gate_46(G575,G5);
not gate_47(G1178,G2236);
not gate_48(G1186,G2253);
not gate_49(G1192,G2256);
buf gate_50(G1198,G38);
buf gate_51(G1205,G15);
nand gate_52(G1206,G12,G9);
nand gate_53(G1207,G12,G9);
buf gate_54(G1210,G38);
not gate_55(G1458,G1455);
not gate_56(G1461,G1459);
buf gate_57(G436,G1462);
not gate_58(G1464,G1462);
not gate_59(G1471,G1469);
buf gate_60(G1475,G106);
not gate_61(G1482,G1480);
not gate_62(G1488,G1486);
not gate_63(G1495,G1492);
not gate_64(G1499,G1496);
not gate_65(G1500,G106);
buf gate_66(G1503,G18);
buf gate_67(G1512,G18);
and gate_68(G1518,G4528,G1492);
buf gate_69(G1524,G18);
not gate_70(G1535,G18);
nand gate_71(G1541,G4528,G1496);
not gate_72(G2207,G2204);
not gate_73(G2210,G2208);
buf gate_74(G478,G2211);
not gate_75(G2213,G2211);
not gate_76(G2220,G2218);
not gate_77(G2226,G2224);
not gate_78(G2232,G2230);
not gate_79(G2238,G2236);
not gate_80(G2241,G2239);
not gate_81(G2249,G2247);
not gate_82(G2255,G2253);
not gate_83(G2258,G2256);
buf gate_84(G2828,G4526);
not gate_85(G3700,G3698);
not gate_86(G3703,G3701);
not gate_87(G3707,G3705);
not gate_88(G3713,G3711);
not gate_89(G3719,G3717);
not gate_90(G3725,G3723);
not gate_91(G3731,G3729);
not gate_92(G3739,G3737);
not gate_93(G3745,G3743);
not gate_94(G3751,G3749);
not gate_95(G4121,G4393);
buf gate_96(G522,G4394);
not gate_97(G4396,G4394);
not gate_98(G4402,G4400);
not gate_99(G4407,G4405);
not gate_100(G4412,G4410);
not gate_101(G4417,G4415);
not gate_102(G4422,G4420);
not gate_103(G4429,G4427);
not gate_104(G4434,G4432);
not gate_105(G4439,G4437);
buf gate_106(G4833,G4526);
nand gate_107(G402,G400,G401);
not gate_108(G404,G2857);
not gate_109(G406,G4514);
not gate_110(G408,G4442);
not gate_111(G410,G1501);
and gate_112(G2876,G2857,G4514);
and gate_113(G2878,G4442,G1501);
buf gate_114(G432,G573);
buf gate_115(G446,G1475);
not gate_116(G1519,G1518);
and gate_117(G2871,G4528,G1458);
nand gate_118(G2883,G4528,G2207);
and gate_119(G280,G1184,G575);
nand gate_120(G284,G1197,G574);
not gate_121(G286,G1205);
nand gate_122(G289,G1197,G574);
nand gate_123(G292,G1184,G575);
not gate_124(G341,G1205);
not gate_125(G4839,G4833);
buf gate_126(G572,G573);
buf gate_127(G581,G1206);
buf gate_128(G587,G1512);
buf gate_129(G601,G1206);
buf gate_130(G606,G1512);
buf gate_131(G650,G1206);
buf gate_132(G657,G1512);
buf gate_133(G671,G1207);
buf gate_134(G678,G1503);
and gate_135(G777,G1541,G1198);
and gate_136(G1115,G1541,G1198);
buf gate_137(G1336,G1512);
buf gate_138(G1350,G1503);
not gate_139(G1477,G1475);
not gate_140(G1507,G1503);
not gate_141(G1514,G1512);
not gate_142(G1530,G1524);
buf gate_143(G2259,G1535);
not gate_144(G2833,G2828);
not gate_145(G2872,G2871);
buf gate_146(G2886,G1207);
buf gate_147(G2892,G1503);
buf gate_148(G2905,G1207);
buf gate_149(G2909,G1503);
buf gate_150(G3622,G1524);
buf gate_151(G3635,G1524);
buf gate_152(G3755,G1535);
buf gate_153(G4640,G1524);
buf gate_154(G4653,G1524);
buf gate_155(G4873,G1541);
buf gate_156(G4876,G1198);
buf gate_157(G4881,G1488);
buf gate_158(G4889,G1482);
buf gate_159(G4905,G1471);
buf gate_160(G4916,G1198);
buf gate_161(G4921,G1464);
buf gate_162(G5175,G1541);
buf gate_163(G5178,G1198);
buf gate_164(G5186,G1198);
buf gate_165(G5191,G1488);
buf gate_166(G5199,G1482);
buf gate_167(G5215,G1471);
buf gate_168(G5223,G1464);
buf gate_169(G5393,G1192);
buf gate_170(G5401,G1186);
buf gate_171(G5409,G2249);
buf gate_172(G5417,G1178);
buf gate_173(G5425,G2232);
buf gate_174(G5433,G2226);
buf gate_175(G5441,G2220);
buf gate_176(G5449,G2241);
buf gate_177(G5457,G2213);
buf gate_178(G5745,G1192);
buf gate_179(G5753,G1186);
buf gate_180(G5761,G2249);
buf gate_181(G5769,G2241);
buf gate_182(G5777,G1178);
buf gate_183(G5785,G2232);
buf gate_184(G5793,G2226);
buf gate_185(G5801,G2220);
buf gate_186(G5809,G2213);
buf gate_187(G5865,G3751);
buf gate_188(G5873,G3745);
buf gate_189(G5881,G3739);
buf gate_190(G5889,G3731);
buf gate_191(G5897,G3725);
buf gate_192(G5905,G3719);
buf gate_193(G5913,G3713);
buf gate_194(G5921,G3707);
buf gate_195(G5985,G3751);
buf gate_196(G5993,G3745);
buf gate_197(G6001,G3739);
buf gate_198(G6009,G3725);
buf gate_199(G6017,G3719);
buf gate_200(G6025,G3713);
buf gate_201(G6033,G3707);
buf gate_202(G6041,G3731);
buf gate_203(G6514,G1210);
buf gate_204(G6554,G1210);
buf gate_205(G6567,G4439);
buf gate_206(G6575,G4434);
buf gate_207(G6583,G4429);
buf gate_208(G6591,G4422);
buf gate_209(G6599,G4417);
buf gate_210(G6607,G4412);
buf gate_211(G6615,G4407);
buf gate_212(G6623,G4402);
buf gate_213(G6631,G4396);
buf gate_214(G6853,G4439);
buf gate_215(G6861,G4434);
buf gate_216(G6869,G4429);
buf gate_217(G6877,G4417);
buf gate_218(G6885,G4412);
buf gate_219(G6893,G4407);
buf gate_220(G6901,G4402);
buf gate_221(G6909,G4422);
buf gate_222(G6917,G4396);
not gate_223(G281,G280);
buf gate_224(G453,G572);
and gate_225(G784,G1519,G1198);
and gate_226(G1014,G1198,G1519);
and gate_227(G3221,G2883,G1210);
buf gate_228(G4913,G1519);
nor gate_229(G4929,G1519,G1198);
buf gate_230(G5183,G1519);
nor gate_231(G5231,G1198,G1519);
buf gate_232(G6511,G2883);
and gate_233(G278,G163,G572);
and gate_234(G615,G170,G587);
not gate_235(G594,G587);
not gate_236(G611,G606);
and gate_237(G617,G169,G587);
and gate_238(G619,G168,G587);
and gate_239(G621,G167,G587);
and gate_240(G623,G166,G606);
and gate_241(G625,G165,G606);
and gate_242(G627,G164,G606);
not gate_243(G664,G657);
not gate_244(G685,G678);
and gate_245(G691,G177,G657);
and gate_246(G693,G176,G657);
and gate_247(G695,G175,G657);
and gate_248(G697,G174,G657);
and gate_249(G699,G173,G657);
and gate_250(G701,G157,G678);
and gate_251(G703,G156,G678);
and gate_252(G705,G155,G678);
and gate_253(G707,G154,G678);
and gate_254(G709,G153,G678);
not gate_255(G4879,G4873);
not gate_256(G4880,G4876);
not gate_257(G4887,G4881);
not gate_258(G4895,G4889);
not gate_259(G4911,G4905);
not gate_260(G4920,G4916);
not gate_261(G4927,G4921);
not gate_262(G5181,G5175);
not gate_263(G5182,G5178);
not gate_264(G5190,G5186);
not gate_265(G5197,G5191);
not gate_266(G5205,G5199);
not gate_267(G5221,G5215);
not gate_268(G5229,G5223);
not gate_269(G1343,G1336);
not gate_270(G1357,G1350);
and gate_271(G1364,G181,G1336);
and gate_272(G1366,G171,G1336);
and gate_273(G1368,G180,G1336);
and gate_274(G1370,G179,G1336);
and gate_275(G1372,G178,G1336);
and gate_276(G1374,G161,G1350);
and gate_277(G1376,G151,G1350);
and gate_278(G1378,G160,G1350);
and gate_279(G1380,G159,G1350);
and gate_280(G1382,G158,G1350);
not gate_281(G5399,G5393);
not gate_282(G5407,G5401);
not gate_283(G5415,G5409);
not gate_284(G5423,G5417);
not gate_285(G5431,G5425);
not gate_286(G5439,G5433);
not gate_287(G5447,G5441);
not gate_288(G5455,G5449);
not gate_289(G5463,G5457);
not gate_290(G5751,G5745);
not gate_291(G5759,G5753);
not gate_292(G5767,G5761);
not gate_293(G5775,G5769);
not gate_294(G5783,G5777);
not gate_295(G5791,G5785);
not gate_296(G5799,G5793);
not gate_297(G5807,G5801);
not gate_298(G5815,G5809);
buf gate_299(G2019,G1514);
buf gate_300(G2032,G1507);
buf gate_301(G2117,G1514);
buf gate_302(G2130,G1507);
not gate_303(G2266,G2259);
buf gate_304(G2272,G1507);
and gate_305(G2286,G44,G2259);
and gate_306(G2288,G41,G2259);
and gate_307(G2290,G29,G2259);
and gate_308(G2292,G26,G2259);
and gate_309(G2294,G23,G2259);
not gate_310(G5871,G5865);
not gate_311(G5879,G5873);
not gate_312(G5887,G5881);
not gate_313(G5895,G5889);
not gate_314(G5903,G5897);
not gate_315(G5911,G5905);
not gate_316(G5919,G5913);
not gate_317(G5927,G5921);
not gate_318(G5991,G5985);
not gate_319(G5999,G5993);
not gate_320(G6007,G6001);
not gate_321(G6015,G6009);
not gate_322(G6023,G6017);
not gate_323(G6031,G6025);
not gate_324(G6039,G6033);
not gate_325(G6047,G6041);
not gate_326(G2899,G2892);
not gate_327(G2914,G2909);
and gate_328(G2919,G209,G2892);
and gate_329(G2921,G216,G2892);
and gate_330(G2923,G215,G2892);
and gate_331(G2925,G214,G2892);
and gate_332(G2927,G213,G2909);
and gate_333(G2929,G212,G2909);
and gate_334(G2931,G211,G2909);
not gate_335(G6518,G6514);
and gate_336(G3173,G2872,G1210);
not gate_337(G6558,G6554);
not gate_338(G6573,G6567);
not gate_339(G6581,G6575);
not gate_340(G6589,G6583);
not gate_341(G6597,G6591);
not gate_342(G6605,G6599);
not gate_343(G6613,G6607);
not gate_344(G6621,G6615);
not gate_345(G6629,G6623);
not gate_346(G6637,G6631);
not gate_347(G3629,G3622);
not gate_348(G3642,G3635);
and gate_349(G3649,G1461,G3622);
and gate_350(G3651,G1464,G3622);
and gate_351(G3653,G1471,G3622);
and gate_352(G3655,G1500,G3622);
and gate_353(G3657,G1482,G3622);
and gate_354(G3659,G1488,G3635);
and gate_355(G3661,G1495,G3635);
and gate_356(G3663,G1499,G3635);
not gate_357(G3762,G3755);
buf gate_358(G3768,G1507);
and gate_359(G3782,G47,G3755);
and gate_360(G3784,G35,G3755);
and gate_361(G3786,G32,G3755);
and gate_362(G3788,G50,G3755);
and gate_363(G3790,G66,G3755);
not gate_364(G6859,G6853);
not gate_365(G6867,G6861);
not gate_366(G6875,G6869);
not gate_367(G6883,G6877);
not gate_368(G6891,G6885);
not gate_369(G6899,G6893);
not gate_370(G6907,G6901);
not gate_371(G6915,G6909);
not gate_372(G6923,G6917);
buf gate_373(G4094,G1530);
buf gate_374(G4107,G1530);
buf gate_375(G4444,G1530);
buf gate_376(G4457,G1530);
not gate_377(G4647,G4640);
not gate_378(G4660,G4653);
and gate_379(G4667,G2210,G4640);
and gate_380(G4669,G2213,G4640);
and gate_381(G4671,G2220,G4640);
and gate_382(G4673,G2226,G4640);
and gate_383(G4675,G2232,G4640);
and gate_384(G4677,G2238,G4653);
and gate_385(G4679,G2241,G4653);
and gate_386(G4681,G2249,G4653);
and gate_387(G4683,G2255,G4653);
and gate_388(G4685,G2258,G4653);
buf gate_389(G4897,G1477);
buf gate_390(G5207,G1477);
buf gate_391(G6551,G2872);
nand gate_392(G763,G4876,G4879);
nand gate_393(G764,G4873,G4880);
not gate_394(G4919,G4913);
nand gate_395(G886,G4913,G4920);
nand gate_396(G1005,G5178,G5181);
nand gate_397(G1006,G5175,G5182);
not gate_398(G5189,G5183);
nand gate_399(G1018,G5183,G5190);
not gate_400(G5237,G5231);
not gate_401(G6517,G6511);
nand gate_402(G3169,G6511,G6518);
not gate_403(G4935,G4929);
buf gate_404(G4970,G784);
buf gate_405(G5239,G1014);
or gate_406(G577,G594,G615);
or gate_407(G616,G594,G587);
or gate_408(G618,G594,G617);
or gate_409(G620,G594,G619);
or gate_410(G622,G594,G621);
or gate_411(G624,G611,G623);
or gate_412(G626,G611,G625);
or gate_413(G628,G611,G627);
or gate_414(G692,G664,G691);
or gate_415(G694,G664,G693);
or gate_416(G696,G664,G695);
or gate_417(G698,G664,G697);
or gate_418(G700,G664,G699);
or gate_419(G702,G685,G701);
or gate_420(G704,G685,G703);
or gate_421(G706,G685,G705);
or gate_422(G708,G685,G707);
or gate_423(G710,G685,G709);
nand gate_424(G765,G763,G764);
not gate_425(G4903,G4897);
nand gate_426(G885,G4916,G4919);
nand gate_427(G1007,G1005,G1006);
nand gate_428(G1017,G5186,G5189);
not gate_429(G5213,G5207);
and gate_430(G1363,G141,G1343);
and gate_431(G1365,G147,G1343);
and gate_432(G1367,G138,G1343);
and gate_433(G1369,G144,G1343);
and gate_434(G1371,G135,G1343);
and gate_435(G1373,G141,G1357);
and gate_436(G1375,G147,G1357);
and gate_437(G1377,G138,G1357);
and gate_438(G1379,G144,G1357);
and gate_439(G1381,G135,G1357);
not gate_440(G2026,G2019);
not gate_441(G2039,G2032);
and gate_442(G2046,G103,G2019);
and gate_443(G2048,G130,G2019);
and gate_444(G2050,G127,G2019);
and gate_445(G2052,G124,G2019);
and gate_446(G2054,G100,G2019);
and gate_447(G2056,G103,G2032);
and gate_448(G2058,G130,G2032);
and gate_449(G2060,G127,G2032);
and gate_450(G2062,G124,G2032);
and gate_451(G2064,G100,G2032);
not gate_452(G2124,G2117);
not gate_453(G2137,G2130);
and gate_454(G2144,G115,G2117);
and gate_455(G2146,G118,G2117);
and gate_456(G2148,G97,G2117);
and gate_457(G2150,G94,G2117);
and gate_458(G2152,G121,G2117);
and gate_459(G2154,G115,G2130);
and gate_460(G2156,G118,G2130);
and gate_461(G2158,G97,G2130);
and gate_462(G2160,G94,G2130);
and gate_463(G2162,G121,G2130);
not gate_464(G2279,G2272);
and gate_465(G2285,G208,G2266);
and gate_466(G2287,G198,G2266);
and gate_467(G2289,G207,G2266);
and gate_468(G2291,G206,G2266);
and gate_469(G2293,G205,G2266);
and gate_470(G2296,G44,G2272);
and gate_471(G2298,G41,G2272);
and gate_472(G2300,G29,G2272);
and gate_473(G2302,G26,G2272);
and gate_474(G2304,G23,G2272);
or gate_475(G2918,G2899,G2892);
or gate_476(G2920,G2899,G2919);
or gate_477(G2922,G2899,G2921);
or gate_478(G2924,G2899,G2923);
or gate_479(G2926,G2899,G2925);
or gate_480(G2928,G2914,G2927);
or gate_481(G2930,G2914,G2929);
or gate_482(G2932,G2914,G2931);
nand gate_483(G3168,G6514,G6517);
not gate_484(G6557,G6551);
nand gate_485(G3211,G6551,G6558);
and gate_486(G3648,G114,G3629);
and gate_487(G3650,G113,G3629);
and gate_488(G3652,G111,G3629);
and gate_489(G3654,G87,G3629);
and gate_490(G3656,G112,G3629);
and gate_491(G3658,G88,G3642);
and gate_492(G3660,G1455,G3642);
and gate_493(G3662,G2204,G3642);
and gate_494(G3665,G3703,G3642);
and gate_495(G3666,G70,G3642);
not gate_496(G3775,G3768);
and gate_497(G3781,G193,G3762);
and gate_498(G3783,G192,G3762);
and gate_499(G3785,G191,G3762);
and gate_500(G3787,G190,G3762);
and gate_501(G3789,G189,G3762);
and gate_502(G3792,G47,G3768);
and gate_503(G3794,G35,G3768);
and gate_504(G3796,G32,G3768);
and gate_505(G3798,G50,G3768);
and gate_506(G3800,G66,G3768);
not gate_507(G4101,G4094);
not gate_508(G4114,G4107);
and gate_509(G4123,G58,G4094);
and gate_510(G4126,G77,G4094);
and gate_511(G4129,G78,G4094);
and gate_512(G4132,G59,G4094);
and gate_513(G4135,G81,G4094);
and gate_514(G4138,G80,G4107);
and gate_515(G4141,G79,G4107);
and gate_516(G4144,G60,G4107);
and gate_517(G4147,G61,G4107);
and gate_518(G4150,G62,G4107);
not gate_519(G4451,G4444);
not gate_520(G4464,G4457);
and gate_521(G4471,G69,G4444);
and gate_522(G4473,G70,G4444);
and gate_523(G4475,G74,G4444);
and gate_524(G4477,G76,G4444);
and gate_525(G4479,G75,G4444);
and gate_526(G4481,G73,G4457);
and gate_527(G4483,G53,G4457);
and gate_528(G4485,G54,G4457);
and gate_529(G4487,G55,G4457);
and gate_530(G4489,G56,G4457);
and gate_531(G4666,G82,G4647);
and gate_532(G4668,G65,G4647);
and gate_533(G4670,G83,G4647);
and gate_534(G4672,G84,G4647);
and gate_535(G4674,G85,G4647);
and gate_536(G4676,G64,G4660);
and gate_537(G4678,G63,G4660);
and gate_538(G4680,G86,G4660);
and gate_539(G4682,G109,G4660);
and gate_540(G4684,G110,G4660);
and gate_541(G579,G577,G581);
and gate_542(G629,G616,G581);
and gate_543(G633,G618,G581);
and gate_544(G637,G620,G581);
and gate_545(G641,G622,G581);
and gate_546(G645,G624,G601);
and gate_547(G711,G692,G650);
and gate_548(G715,G694,G650);
and gate_549(G719,G696,G650);
and gate_550(G723,G698,G650);
and gate_551(G727,G700,G650);
and gate_552(G731,G702,G671);
and gate_553(G737,G704,G671);
and gate_554(G745,G706,G671);
and gate_555(G751,G708,G671);
and gate_556(G757,G710,G671);
nand gate_557(G887,G885,G886);
nand gate_558(G1019,G1017,G1018);
not gate_559(G5245,G5239);
or gate_560(G1383,G1365,G1366);
or gate_561(G1387,G1367,G1368);
or gate_562(G1391,G1369,G1370);
or gate_563(G1395,G1371,G1372);
or gate_564(G1399,G1375,G1376);
or gate_565(G1406,G1377,G1378);
or gate_566(G1412,G1379,G1380);
or gate_567(G1418,G1381,G1382);
or gate_568(G2305,G2287,G2288);
or gate_569(G2308,G2289,G2290);
or gate_570(G2312,G2291,G2292);
or gate_571(G2316,G2293,G2294);
and gate_572(G2933,G2920,G2886);
and gate_573(G2938,G2922,G2886);
and gate_574(G2942,G2924,G2886);
and gate_575(G2946,G2926,G2886);
and gate_576(G2950,G2928,G2905);
nand gate_577(G3170,G3168,G3169);
nand gate_578(G3210,G6554,G6557);
or gate_579(G3667,G3650,G3651);
or gate_580(G3670,G3652,G3653);
or gate_581(G3673,G3654,G3655);
or gate_582(G3676,G3656,G3657);
or gate_583(G3679,G3658,G3659);
or gate_584(G3682,G3665,G3635);
or gate_585(G3686,G3666,G3635);
or gate_586(G3801,G3781,G3782);
or gate_587(G3804,G3783,G3784);
or gate_588(G3807,G3785,G3786);
or gate_589(G3810,G3787,G3788);
or gate_590(G3813,G3789,G3790);
and gate_591(G4525,G2918,G2886);
or gate_592(G4686,G4668,G4669);
or gate_593(G4689,G4670,G4671);
or gate_594(G4692,G4672,G4673);
or gate_595(G4695,G4674,G4675);
or gate_596(G4698,G4676,G4677);
or gate_597(G4701,G4678,G4679);
or gate_598(G4704,G4680,G4681);
or gate_599(G4707,G4682,G4683);
or gate_600(G4710,G4684,G4685);
not gate_601(G4976,G4970);
and gate_602(G5271,G2932,G2905);
and gate_603(G5274,G2930,G2905);
and gate_604(G5305,G628,G601);
and gate_605(G5308,G626,G601);
or gate_606(G5318,G1373,G1374);
or gate_607(G6690,G3648,G3649);
or gate_608(G6711,G3662,G3663);
or gate_609(G6714,G3660,G3661);
or gate_610(G7252,G2285,G2286);
or gate_611(G7296,G1363,G1364);
or gate_612(G7466,G4666,G4667);
and gate_613(G907,G765,G784);
and gate_614(G913,G765,G784);
and gate_615(G915,G765,G784);
and gate_616(G916,G765,G784);
and gate_617(G1116,G1007,G1014);
and gate_618(G2045,G204,G2026);
and gate_619(G2047,G203,G2026);
and gate_620(G2049,G202,G2026);
and gate_621(G2051,G201,G2026);
and gate_622(G2053,G200,G2026);
and gate_623(G2055,G235,G2039);
and gate_624(G2057,G234,G2039);
and gate_625(G2059,G233,G2039);
and gate_626(G2061,G232,G2039);
and gate_627(G2063,G231,G2039);
and gate_628(G2143,G197,G2124);
and gate_629(G2145,G187,G2124);
and gate_630(G2147,G196,G2124);
and gate_631(G2149,G195,G2124);
and gate_632(G2151,G194,G2124);
and gate_633(G2153,G227,G2137);
and gate_634(G2155,G217,G2137);
and gate_635(G2157,G226,G2137);
and gate_636(G2159,G225,G2137);
and gate_637(G2161,G224,G2137);
and gate_638(G2295,G239,G2279);
and gate_639(G2297,G229,G2279);
and gate_640(G2299,G238,G2279);
and gate_641(G2301,G237,G2279);
and gate_642(G2303,G236,G2279);
nand gate_643(G3212,G3210,G3211);
and gate_644(G3791,G223,G3775);
and gate_645(G3793,G222,G3775);
and gate_646(G3795,G221,G3775);
and gate_647(G3797,G220,G3775);
and gate_648(G3799,G219,G3775);
and gate_649(G4122,G4121,G4101);
and gate_650(G4125,G4396,G4101);
and gate_651(G4128,G4402,G4101);
and gate_652(G4131,G4407,G4101);
and gate_653(G4134,G4412,G4101);
and gate_654(G4137,G4417,G4114);
and gate_655(G4140,G4422,G4114);
and gate_656(G4143,G4429,G4114);
and gate_657(G4146,G4434,G4114);
and gate_658(G4149,G4439,G4114);
and gate_659(G4470,G3700,G4451);
and gate_660(G4472,G3703,G4451);
and gate_661(G4474,G3707,G4451);
and gate_662(G4476,G3713,G4451);
and gate_663(G4478,G3719,G4451);
and gate_664(G4480,G3725,G4464);
and gate_665(G4482,G3731,G4464);
and gate_666(G4484,G3739,G4464);
and gate_667(G4486,G3745,G4464);
and gate_668(G4488,G3751,G4464);
buf gate_669(G4962,G765);
buf gate_670(G5003,G765);
buf gate_671(G5234,G1007);
buf gate_672(G5242,G1007);
not gate_673(G5250,G4525);
not gate_674(G5284,G579);
and gate_675(G802,G1488,G2950);
and gate_676(G821,G1482,G2946);
and gate_677(G845,G1477,G2942);
and gate_678(G868,G1471,G2938);
and gate_679(G877,G1464,G2933);
and gate_680(G902,G887,G765);
or gate_681(G908,G777,G907);
and gate_682(G914,G887,G765);
or gate_683(G917,G777,G916);
and gate_684(G953,G887,G765);
not gate_685(G1023,G1019);
and gate_686(G1035,G1488,G2950);
and gate_687(G1050,G1482,G2946);
and gate_688(G1068,G1477,G2942);
and gate_689(G1086,G1471,G2938);
and gate_690(G1102,G1464,G2933);
and gate_691(G1108,G1019,G1007);
or gate_692(G1117,G1115,G1116);
not gate_693(G5322,G5318);
and gate_694(G1553,G1192,G757);
and gate_695(G1567,G1186,G751);
and gate_696(G1584,G2249,G745);
and gate_697(G1590,G2241,G737);
and gate_698(G1606,G1178,G731);
and gate_699(G1624,G2232,G1418);
and gate_700(G1647,G2226,G1412);
and gate_701(G1669,G2220,G1406);
and gate_702(G1677,G2213,G1399);
and gate_703(G1802,G1192,G757);
and gate_704(G1816,G1186,G751);
and gate_705(G1834,G2249,G745);
and gate_706(G1841,G737,G2241);
and gate_707(G1866,G1178,G731);
and gate_708(G1880,G2232,G1418);
and gate_709(G1897,G2226,G1412);
and gate_710(G1914,G2220,G1406);
and gate_711(G1929,G2213,G1399);
or gate_712(G2065,G2045,G2046);
or gate_713(G2069,G2047,G2048);
or gate_714(G2073,G2049,G2050);
or gate_715(G2077,G2051,G2052);
or gate_716(G2081,G2053,G2054);
or gate_717(G2085,G2055,G2056);
or gate_718(G2091,G2057,G2058);
or gate_719(G2099,G2059,G2060);
or gate_720(G2105,G2061,G2062);
or gate_721(G2111,G2063,G2064);
or gate_722(G2163,G2145,G2146);
or gate_723(G2167,G2147,G2148);
or gate_724(G2171,G2149,G2150);
or gate_725(G2175,G2151,G2152);
or gate_726(G2179,G2155,G2156);
or gate_727(G2186,G2157,G2158);
or gate_728(G2192,G2159,G2160);
or gate_729(G2198,G2161,G2162);
or gate_730(G2320,G2297,G2298);
or gate_731(G2323,G2299,G2300);
or gate_732(G2329,G2301,G2302);
or gate_733(G2335,G2303,G2304);
and gate_734(G2962,G4710,G727);
and gate_735(G2970,G4707,G723);
and gate_736(G2977,G4704,G719);
and gate_737(G2979,G4701,G715);
and gate_738(G2989,G4698,G711);
and gate_739(G2998,G4695,G1395);
and gate_740(G3006,G4692,G1391);
and gate_741(G3013,G4689,G1387);
and gate_742(G3015,G4686,G1383);
and gate_743(G3183,G3679,G645);
and gate_744(G3192,G3676,G641);
and gate_745(G3200,G3673,G637);
and gate_746(G3207,G3670,G633);
and gate_747(G3209,G3667,G629);
and gate_748(G3216,G3212,G3170);
and gate_749(G3222,G3170,G3173);
not gate_750(G6694,G6690);
and gate_751(G3695,G1535,G2305);
or gate_752(G3816,G3791,G3792);
or gate_753(G3821,G3793,G3794);
or gate_754(G3828,G3795,G3796);
or gate_755(G3833,G3797,G3798);
or gate_756(G3838,G3799,G3800);
or gate_757(G4151,G4125,G4126);
or gate_758(G4154,G4128,G4129);
or gate_759(G4157,G4131,G4132);
or gate_760(G4160,G4134,G4135);
or gate_761(G4163,G4137,G4138);
or gate_762(G4166,G4140,G4141);
or gate_763(G4169,G4143,G4144);
or gate_764(G4172,G4146,G4147);
or gate_765(G4175,G4149,G4150);
not gate_766(G7256,G7252);
not gate_767(G7300,G7296);
or gate_768(G4490,G4474,G4475);
or gate_769(G4493,G4476,G4477);
or gate_770(G4496,G4478,G4479);
or gate_771(G4499,G4480,G4481);
or gate_772(G4502,G4482,G4483);
or gate_773(G4505,G4484,G4485);
or gate_774(G4508,G4486,G4487);
or gate_775(G4511,G4488,G4489);
not gate_776(G7470,G7466);
buf gate_777(G4884,G2950);
buf gate_778(G4892,G2946);
buf gate_779(G4900,G2942);
buf gate_780(G4908,G2938);
buf gate_781(G4924,G2933);
buf gate_782(G4952,G887);
nor gate_783(G4983,G777,G915);
buf gate_784(G4993,G887);
nor gate_785(G5011,G1464,G2933);
buf gate_786(G5194,G2950);
buf gate_787(G5202,G2946);
buf gate_788(G5210,G2942);
buf gate_789(G5218,G2938);
buf gate_790(G5226,G2933);
buf gate_791(G5247,G2933);
buf gate_792(G5255,G2942);
buf gate_793(G5258,G2938);
buf gate_794(G5263,G2950);
buf gate_795(G5266,G2946);
not gate_796(G5277,G5271);
not gate_797(G5278,G5274);
buf gate_798(G5281,G629);
buf gate_799(G5289,G637);
buf gate_800(G5292,G633);
buf gate_801(G5297,G645);
buf gate_802(G5300,G641);
not gate_803(G5311,G5305);
not gate_804(G5312,G5308);
buf gate_805(G5315,G1399);
buf gate_806(G5323,G1412);
buf gate_807(G5326,G1406);
buf gate_808(G5331,G731);
buf gate_809(G5334,G1418);
buf gate_810(G5339,G745);
buf gate_811(G5342,G737);
buf gate_812(G5349,G757);
buf gate_813(G5352,G751);
buf gate_814(G5396,G757);
buf gate_815(G5404,G751);
buf gate_816(G5412,G745);
buf gate_817(G5420,G731);
buf gate_818(G5428,G1418);
buf gate_819(G5436,G1412);
buf gate_820(G5444,G1406);
buf gate_821(G5452,G737);
buf gate_822(G5460,G1399);
nor gate_823(G5465,G2241,G737);
nor gate_824(G5581,G2213,G1399);
buf gate_825(G5748,G757);
buf gate_826(G5756,G751);
buf gate_827(G5764,G745);
buf gate_828(G5772,G737);
buf gate_829(G5780,G731);
buf gate_830(G5788,G1418);
buf gate_831(G5796,G1412);
buf gate_832(G5804,G1406);
buf gate_833(G5812,G1399);
nor gate_834(G5849,G737,G2241);
buf gate_835(G5929,G3682);
buf gate_836(G6049,G3682);
buf gate_837(G6367,G4710);
buf gate_838(G6370,G727);
buf gate_839(G6375,G4707);
buf gate_840(G6378,G723);
buf gate_841(G6383,G4704);
buf gate_842(G6386,G719);
buf gate_843(G6391,G4698);
buf gate_844(G6394,G711);
buf gate_845(G6399,G4695);
buf gate_846(G6402,G1395);
buf gate_847(G6407,G4692);
buf gate_848(G6410,G1391);
buf gate_849(G6415,G4689);
buf gate_850(G6418,G1387);
buf gate_851(G6423,G4701);
buf gate_852(G6426,G715);
buf gate_853(G6431,G4686);
buf gate_854(G6434,G1383);
buf gate_855(G6442,G3813);
buf gate_856(G6450,G3810);
buf gate_857(G6458,G3807);
buf gate_858(G6466,G3801);
buf gate_859(G6498,G3804);
buf gate_860(G6519,G3679);
buf gate_861(G6522,G645);
buf gate_862(G6527,G3676);
buf gate_863(G6530,G641);
buf gate_864(G6535,G3673);
buf gate_865(G6538,G637);
buf gate_866(G6543,G3670);
buf gate_867(G6546,G633);
buf gate_868(G6559,G3667);
buf gate_869(G6562,G629);
buf gate_870(G6687,G3667);
buf gate_871(G6695,G3673);
buf gate_872(G6698,G3670);
buf gate_873(G6703,G3679);
buf gate_874(G6706,G3676);
not gate_875(G6717,G6711);
not gate_876(G6718,G6714);
or gate_877(G6724,G2153,G2154);
or gate_878(G6768,G2295,G2296);
or gate_879(G7208,G2143,G2144);
buf gate_880(G7221,G3801);
buf gate_881(G7229,G3807);
buf gate_882(G7232,G3804);
buf gate_883(G7239,G3813);
buf gate_884(G7242,G3810);
buf gate_885(G7249,G2305);
buf gate_886(G7257,G2312);
buf gate_887(G7260,G2308);
buf gate_888(G7268,G2316);
buf gate_889(G7293,G1383);
buf gate_890(G7301,G1391);
buf gate_891(G7304,G1387);
buf gate_892(G7309,G711);
buf gate_893(G7312,G1395);
buf gate_894(G7317,G719);
buf gate_895(G7320,G715);
buf gate_896(G7327,G727);
buf gate_897(G7330,G723);
buf gate_898(G7396,G2316);
buf gate_899(G7404,G2312);
buf gate_900(G7412,G2308);
buf gate_901(G7425,G3686);
buf gate_902(G7463,G4686);
buf gate_903(G7471,G4692);
buf gate_904(G7474,G4689);
buf gate_905(G7479,G4698);
buf gate_906(G7482,G4695);
buf gate_907(G7487,G4704);
buf gate_908(G7490,G4701);
buf gate_909(G7497,G4710);
buf gate_910(G7500,G4707);
or gate_911(G7507,G4472,G4473);
or gate_912(G7510,G4470,G4471);
or gate_913(G7554,G4122,G4123);
nand gate_914(G1152,G5234,G5237);
not gate_915(G5238,G5234);
nand gate_916(G1156,G5242,G5245);
not gate_917(G5246,G5242);
not gate_918(G5254,G5250);
not gate_919(G5288,G5284);
or gate_920(G3223,G3221,G3222);
or gate_921(G4942,G777,G913,G914);
not gate_922(G4966,G4962);
not gate_923(G5007,G5003);
nand gate_924(G5279,G5274,G5277);
nand gate_925(G5280,G5271,G5278);
nand gate_926(G5313,G5308,G5311);
nand gate_927(G5314,G5305,G5312);
nand gate_928(G6719,G6714,G6717);
nand gate_929(G6720,G6711,G6718);
nand gate_930(G790,G4884,G4887);
not gate_931(G4888,G4884);
nand gate_932(G803,G4892,G4895);
not gate_933(G4896,G4892);
nand gate_934(G825,G4900,G4903);
not gate_935(G4904,G4900);
nand gate_936(G851,G4908,G4911);
not gate_937(G4912,G4908);
nand gate_938(G893,G4924,G4927);
not gate_939(G4928,G4924);
not gate_940(G906,G902);
not gate_941(G912,G908);
nand gate_942(G1024,G5194,G5197);
not gate_943(G5198,G5194);
nand gate_944(G1036,G5202,G5205);
not gate_945(G5206,G5202);
nand gate_946(G1053,G5210,G5213);
not gate_947(G5214,G5210);
nand gate_948(G1072,G5218,G5221);
not gate_949(G5222,G5218);
nand gate_950(G1091,G5226,G5229);
not gate_951(G5230,G5226);
not gate_952(G1112,G1108);
not gate_953(G1121,G1117);
nand gate_954(G1153,G5231,G5238);
nand gate_955(G1157,G5239,G5246);
not gate_956(G5253,G5247);
nand gate_957(G1216,G5247,G5254);
not gate_958(G5261,G5255);
not gate_959(G5262,G5258);
not gate_960(G5269,G5263);
not gate_961(G5270,G5266);
not gate_962(G5287,G5281);
nand gate_963(G1239,G5281,G5288);
not gate_964(G5295,G5289);
not gate_965(G5296,G5292);
not gate_966(G5303,G5297);
not gate_967(G5304,G5300);
not gate_968(G5321,G5315);
nand gate_969(G1262,G5315,G5322);
not gate_970(G5329,G5323);
not gate_971(G5330,G5326);
not gate_972(G5337,G5331);
not gate_973(G5338,G5334);
nand gate_974(G1544,G5396,G5399);
not gate_975(G5400,G5396);
nand gate_976(G1554,G5404,G5407);
not gate_977(G5408,G5404);
nand gate_978(G1571,G5412,G5415);
not gate_979(G5416,G5412);
nand gate_980(G1596,G5420,G5423);
not gate_981(G5424,G5420);
nand gate_982(G1607,G5428,G5431);
not gate_983(G5432,G5428);
nand gate_984(G1628,G5436,G5439);
not gate_985(G5440,G5436);
nand gate_986(G1653,G5444,G5447);
not gate_987(G5448,G5444);
nand gate_988(G1685,G5452,G5455);
not gate_989(G5456,G5452);
nand gate_990(G1693,G5460,G5463);
not gate_991(G5464,G5460);
nand gate_992(G1793,G5748,G5751);
not gate_993(G5752,G5748);
nand gate_994(G1803,G5756,G5759);
not gate_995(G5760,G5756);
nand gate_996(G1820,G5764,G5767);
not gate_997(G5768,G5764);
nand gate_998(G1848,G5772,G5775);
not gate_999(G5776,G5772);
nand gate_1000(G1857,G5780,G5783);
not gate_1001(G5784,G5780);
nand gate_1002(G1867,G5788,G5791);
not gate_1003(G5792,G5788);
nand gate_1004(G1883,G5796,G5799);
not gate_1005(G5800,G5796);
nand gate_1006(G1901,G5804,G5807);
not gate_1007(G5808,G5804);
nand gate_1008(G1919,G5812,G5815);
not gate_1009(G5816,G5812);
not gate_1010(G5855,G5849);
and gate_1011(G2351,G3751,G2111);
and gate_1012(G2366,G3745,G2105);
and gate_1013(G2384,G3739,G2099);
and gate_1014(G2391,G2091,G3731);
and gate_1015(G2417,G3725,G2085);
and gate_1016(G2431,G3719,G2335);
and gate_1017(G2448,G3713,G2329);
and gate_1018(G2465,G3707,G2323);
not gate_1019(G5935,G5929);
and gate_1020(G2597,G3751,G2111);
and gate_1021(G2612,G3745,G2105);
and gate_1022(G2629,G3739,G2099);
and gate_1023(G2635,G3731,G2091);
and gate_1024(G2652,G3725,G2085);
and gate_1025(G2670,G3719,G2335);
and gate_1026(G2693,G3713,G2329);
and gate_1027(G2715,G3707,G2323);
not gate_1028(G6055,G6049);
not gate_1029(G6373,G6367);
not gate_1030(G6374,G6370);
not gate_1031(G6381,G6375);
not gate_1032(G6382,G6378);
not gate_1033(G6389,G6383);
not gate_1034(G6390,G6386);
not gate_1035(G6397,G6391);
not gate_1036(G6398,G6394);
not gate_1037(G6405,G6399);
not gate_1038(G6406,G6402);
not gate_1039(G6413,G6407);
not gate_1040(G6414,G6410);
not gate_1041(G6421,G6415);
not gate_1042(G6422,G6418);
not gate_1043(G6429,G6423);
not gate_1044(G6430,G6426);
not gate_1045(G6437,G6431);
not gate_1046(G6438,G6434);
not gate_1047(G6446,G6442);
and gate_1048(G3059,G4175,G3813);
not gate_1049(G6454,G6450);
and gate_1050(G3068,G4172,G3810);
not gate_1051(G6462,G6458);
and gate_1052(G3076,G4169,G3807);
and gate_1053(G3079,G4166,G3804);
not gate_1054(G6470,G6466);
and gate_1055(G3090,G4163,G3801);
and gate_1056(G3099,G4160,G2175);
and gate_1057(G3107,G4157,G2171);
and gate_1058(G3114,G4154,G2167);
and gate_1059(G3116,G4151,G2163);
not gate_1060(G6502,G6498);
not gate_1061(G6525,G6519);
not gate_1062(G6526,G6522);
not gate_1063(G6533,G6527);
not gate_1064(G6534,G6530);
not gate_1065(G6541,G6535);
not gate_1066(G6542,G6538);
not gate_1067(G6549,G6543);
not gate_1068(G6550,G6546);
not gate_1069(G6565,G6559);
not gate_1070(G6566,G6562);
not gate_1071(G3220,G3216);
and gate_1072(G3292,G4439,G3838);
and gate_1073(G3308,G4434,G3833);
and gate_1074(G3327,G4429,G3828);
and gate_1075(G3335,G3821,G4422);
and gate_1076(G3362,G4417,G3816);
and gate_1077(G3376,G4412,G2198);
and gate_1078(G3393,G4407,G2192);
and gate_1079(G3410,G4402,G2186);
and gate_1080(G3425,G4396,G2179);
not gate_1081(G6693,G6687);
nand gate_1082(G3503,G6687,G6694);
not gate_1083(G6701,G6695);
not gate_1084(G6702,G6698);
not gate_1085(G6709,G6703);
not gate_1086(G6710,G6706);
not gate_1087(G6728,G6724);
not gate_1088(G6772,G6768);
and gate_1089(G3853,G4439,G3838);
and gate_1090(G3868,G4434,G3833);
and gate_1091(G3885,G4429,G3828);
and gate_1092(G3891,G4422,G3821);
and gate_1093(G3908,G4417,G3816);
and gate_1094(G3926,G4412,G2198);
and gate_1095(G3949,G4407,G2192);
and gate_1096(G3971,G4402,G2186);
and gate_1097(G3979,G4396,G2179);
not gate_1098(G7212,G7208);
not gate_1099(G7227,G7221);
not gate_1100(G7255,G7249);
nand gate_1101(G4202,G7249,G7256);
not gate_1102(G7263,G7257);
not gate_1103(G7264,G7260);
not gate_1104(G7272,G7268);
not gate_1105(G7299,G7293);
nand gate_1106(G4225,G7293,G7300);
not gate_1107(G7307,G7301);
not gate_1108(G7308,G7304);
not gate_1109(G7315,G7309);
not gate_1110(G7316,G7312);
and gate_1111(G4297,G4511,G2081);
and gate_1112(G4305,G4508,G2077);
and gate_1113(G4312,G4505,G2073);
and gate_1114(G4314,G4502,G2069);
and gate_1115(G4324,G4499,G2065);
not gate_1116(G7400,G7396);
and gate_1117(G4333,G4496,G2316);
not gate_1118(G7408,G7404);
and gate_1119(G4341,G4493,G2312);
not gate_1120(G7416,G7412);
and gate_1121(G4348,G4490,G2308);
and gate_1122(G4349,G3686,G3695);
not gate_1123(G7431,G7425);
and gate_1124(G4389,G2320,G1535);
not gate_1125(G7469,G7463);
nand gate_1126(G4530,G7463,G7470);
not gate_1127(G7477,G7471);
not gate_1128(G7478,G7474);
not gate_1129(G7485,G7479);
not gate_1130(G7486,G7482);
not gate_1131(G7513,G7507);
not gate_1132(G7514,G7510);
not gate_1133(G7558,G7554);
or gate_1134(G4932,G917,G953);
not gate_1135(G4956,G4952);
not gate_1136(G4973,G917);
not gate_1137(G4987,G4983);
not gate_1138(G4997,G4993);
not gate_1139(G5017,G5011);
buf gate_1140(G5099,G877);
not gate_1141(G5345,G5339);
not gate_1142(G5346,G5342);
not gate_1143(G5355,G5349);
not gate_1144(G5356,G5352);
nand gate_1145(G5372,G5279,G5280);
nand gate_1146(G5380,G5313,G5314);
not gate_1147(G5471,G5465);
buf gate_1148(G5523,G1590);
not gate_1149(G5587,G5581);
buf gate_1150(G5669,G1677);
buf gate_1151(G5857,G1841);
buf gate_1152(G5868,G2111);
buf gate_1153(G5876,G2105);
buf gate_1154(G5884,G2099);
buf gate_1155(G5892,G2091);
buf gate_1156(G5900,G2085);
buf gate_1157(G5908,G2335);
buf gate_1158(G5916,G2329);
buf gate_1159(G5924,G2323);
nor gate_1160(G5969,G2091,G3731);
buf gate_1161(G5988,G2111);
buf gate_1162(G5996,G2105);
buf gate_1163(G6004,G2099);
buf gate_1164(G6012,G2085);
buf gate_1165(G6020,G2335);
buf gate_1166(G6028,G2329);
buf gate_1167(G6036,G2323);
buf gate_1168(G6044,G2091);
nor gate_1169(G6057,G3731,G2091);
buf gate_1170(G6439,G4175);
buf gate_1171(G6447,G4172);
buf gate_1172(G6455,G4169);
buf gate_1173(G6463,G4163);
buf gate_1174(G6471,G4160);
buf gate_1175(G6474,G2175);
buf gate_1176(G6479,G4157);
buf gate_1177(G6482,G2171);
buf gate_1178(G6487,G4154);
buf gate_1179(G6490,G2167);
buf gate_1180(G6495,G4166);
buf gate_1181(G6503,G4151);
buf gate_1182(G6506,G2163);
buf gate_1183(G6570,G3838);
buf gate_1184(G6578,G3833);
buf gate_1185(G6586,G3828);
buf gate_1186(G6594,G3821);
buf gate_1187(G6602,G3816);
buf gate_1188(G6610,G2198);
buf gate_1189(G6618,G2192);
buf gate_1190(G6626,G2186);
buf gate_1191(G6634,G2179);
nor gate_1192(G6671,G3821,G4422);
buf gate_1193(G6721,G2179);
buf gate_1194(G6729,G2192);
buf gate_1195(G6732,G2186);
buf gate_1196(G6737,G3816);
buf gate_1197(G6740,G2198);
buf gate_1198(G6745,G3828);
buf gate_1199(G6748,G3821);
buf gate_1200(G6755,G3838);
buf gate_1201(G6758,G3833);
buf gate_1202(G6765,G2320);
buf gate_1203(G6773,G2329);
buf gate_1204(G6776,G2323);
buf gate_1205(G6781,G2085);
buf gate_1206(G6784,G2335);
buf gate_1207(G6789,G2099);
buf gate_1208(G6792,G2091);
buf gate_1209(G6799,G2111);
buf gate_1210(G6802,G2105);
nand gate_1211(G6832,G6719,G6720);
buf gate_1212(G6856,G3838);
buf gate_1213(G6864,G3833);
buf gate_1214(G6872,G3828);
buf gate_1215(G6880,G3816);
buf gate_1216(G6888,G2198);
buf gate_1217(G6896,G2192);
buf gate_1218(G6904,G2186);
buf gate_1219(G6912,G3821);
buf gate_1220(G6920,G2179);
nor gate_1221(G6925,G4422,G3821);
nor gate_1222(G7041,G4396,G2179);
buf gate_1223(G7205,G2163);
buf gate_1224(G7213,G2171);
buf gate_1225(G7216,G2167);
buf gate_1226(G7224,G2175);
not gate_1227(G7235,G7229);
not gate_1228(G7236,G7232);
not gate_1229(G7245,G7239);
not gate_1230(G7246,G7242);
buf gate_1231(G7265,G2065);
buf gate_1232(G7273,G2073);
buf gate_1233(G7276,G2069);
buf gate_1234(G7283,G2081);
buf gate_1235(G7286,G2077);
not gate_1236(G7323,G7317);
not gate_1237(G7324,G7320);
not gate_1238(G7333,G7327);
not gate_1239(G7334,G7330);
buf gate_1240(G7361,G4511);
buf gate_1241(G7364,G2081);
buf gate_1242(G7369,G4508);
buf gate_1243(G7372,G2077);
buf gate_1244(G7377,G4505);
buf gate_1245(G7380,G2073);
buf gate_1246(G7385,G4499);
buf gate_1247(G7388,G2065);
buf gate_1248(G7393,G4496);
buf gate_1249(G7401,G4493);
buf gate_1250(G7409,G4490);
buf gate_1251(G7417,G4502);
buf gate_1252(G7420,G2069);
buf gate_1253(G7428,G3695);
not gate_1254(G7493,G7487);
not gate_1255(G7494,G7490);
not gate_1256(G7503,G7497);
not gate_1257(G7504,G7500);
buf gate_1258(G7515,G4493);
buf gate_1259(G7518,G4490);
buf gate_1260(G7523,G4499);
buf gate_1261(G7526,G4496);
buf gate_1262(G7531,G4505);
buf gate_1263(G7534,G4502);
buf gate_1264(G7541,G4511);
buf gate_1265(G7544,G4508);
buf gate_1266(G7551,G4151);
buf gate_1267(G7559,G4157);
buf gate_1268(G7562,G4154);
buf gate_1269(G7567,G4163);
buf gate_1270(G7570,G4160);
buf gate_1271(G7575,G4169);
buf gate_1272(G7578,G4166);
buf gate_1273(G7585,G4175);
buf gate_1274(G7588,G4172);
nand gate_1275(G1176,G1121,G1112);
nand gate_1276(G957,G912,G906);
nand gate_1277(G791,G4881,G4888);
nand gate_1278(G804,G4889,G4896);
nand gate_1279(G826,G4897,G4904);
nand gate_1280(G852,G4905,G4912);
nand gate_1281(G894,G4921,G4928);
nand gate_1282(G1025,G5191,G5198);
nand gate_1283(G1037,G5199,G5206);
nand gate_1284(G1054,G5207,G5214);
nand gate_1285(G1073,G5215,G5222);
nand gate_1286(G1092,G5223,G5230);
nand gate_1287(G1154,G1152,G1153);
nand gate_1288(G1158,G1156,G1157);
nand gate_1289(G1215,G5250,G5253);
nand gate_1290(G1224,G5258,G5261);
nand gate_1291(G1225,G5255,G5262);
nand gate_1292(G1233,G5266,G5269);
nand gate_1293(G1234,G5263,G5270);
nand gate_1294(G1238,G5284,G5287);
nand gate_1295(G1247,G5292,G5295);
nand gate_1296(G1248,G5289,G5296);
nand gate_1297(G1256,G5300,G5303);
nand gate_1298(G1257,G5297,G5304);
nand gate_1299(G1261,G5318,G5321);
nand gate_1300(G1270,G5326,G5329);
nand gate_1301(G1271,G5323,G5330);
nand gate_1302(G1279,G5334,G5337);
nand gate_1303(G1280,G5331,G5338);
nand gate_1304(G1545,G5393,G5400);
nand gate_1305(G1555,G5401,G5408);
nand gate_1306(G1572,G5409,G5416);
nand gate_1307(G1597,G5417,G5424);
nand gate_1308(G1608,G5425,G5432);
nand gate_1309(G1629,G5433,G5440);
nand gate_1310(G1654,G5441,G5448);
nand gate_1311(G1686,G5449,G5456);
nand gate_1312(G1694,G5457,G5464);
nand gate_1313(G1794,G5745,G5752);
nand gate_1314(G1804,G5753,G5760);
nand gate_1315(G1821,G5761,G5768);
nand gate_1316(G1849,G5769,G5776);
nand gate_1317(G1858,G5777,G5784);
nand gate_1318(G1868,G5785,G5792);
nand gate_1319(G1884,G5793,G5800);
nand gate_1320(G1902,G5801,G5808);
nand gate_1321(G1920,G5809,G5816);
nand gate_1322(G2954,G6370,G6373);
nand gate_1323(G2955,G6367,G6374);
nand gate_1324(G2963,G6378,G6381);
nand gate_1325(G2964,G6375,G6382);
nand gate_1326(G2971,G6386,G6389);
nand gate_1327(G2972,G6383,G6390);
nand gate_1328(G2980,G6394,G6397);
nand gate_1329(G2981,G6391,G6398);
nand gate_1330(G2990,G6402,G6405);
nand gate_1331(G2991,G6399,G6406);
nand gate_1332(G2999,G6410,G6413);
nand gate_1333(G3000,G6407,G6414);
nand gate_1334(G3007,G6418,G6421);
nand gate_1335(G3008,G6415,G6422);
nand gate_1336(G3016,G6426,G6429);
nand gate_1337(G3017,G6423,G6430);
nand gate_1338(G3019,G6434,G6437);
nand gate_1339(G3020,G6431,G6438);
nand gate_1340(G3174,G6522,G6525);
nand gate_1341(G3175,G6519,G6526);
nand gate_1342(G3184,G6530,G6533);
nand gate_1343(G3185,G6527,G6534);
nand gate_1344(G3193,G6538,G6541);
nand gate_1345(G3194,G6535,G6542);
nand gate_1346(G3201,G6546,G6549);
nand gate_1347(G3202,G6543,G6550);
nand gate_1348(G3213,G6562,G6565);
nand gate_1349(G3214,G6559,G6566);
not gate_1350(G3227,G3223);
nand gate_1351(G3502,G6690,G6693);
nand gate_1352(G3511,G6698,G6701);
nand gate_1353(G3512,G6695,G6702);
nand gate_1354(G3520,G6706,G6709);
nand gate_1355(G3521,G6703,G6710);
nand gate_1356(G4201,G7252,G7255);
nand gate_1357(G4210,G7260,G7263);
nand gate_1358(G4211,G7257,G7264);
nand gate_1359(G4224,G7296,G7299);
nand gate_1360(G4233,G7304,G7307);
nand gate_1361(G4234,G7301,G7308);
nand gate_1362(G4242,G7312,G7315);
nand gate_1363(G4243,G7309,G7316);
nand gate_1364(G4529,G7466,G7469);
nand gate_1365(G4538,G7474,G7477);
nand gate_1366(G4539,G7471,G7478);
nand gate_1367(G4547,G7482,G7485);
nand gate_1368(G4548,G7479,G7486);
nand gate_1369(G4552,G7510,G7513);
nand gate_1370(G4553,G7507,G7514);
not gate_1371(G4946,G4942);
nand gate_1372(G5347,G5342,G5345);
nand gate_1373(G5348,G5339,G5346);
nand gate_1374(G5357,G5352,G5355);
nand gate_1375(G5358,G5349,G5356);
nand gate_1376(G7237,G7232,G7235);
nand gate_1377(G7238,G7229,G7236);
nand gate_1378(G7247,G7242,G7245);
nand gate_1379(G7248,G7239,G7246);
nand gate_1380(G7325,G7320,G7323);
nand gate_1381(G7326,G7317,G7324);
nand gate_1382(G7335,G7330,G7333);
nand gate_1383(G7336,G7327,G7334);
nand gate_1384(G7495,G7490,G7493);
nand gate_1385(G7496,G7487,G7494);
nand gate_1386(G7505,G7500,G7503);
nand gate_1387(G7506,G7497,G7504);
nand gate_1388(G3244,G3227,G3220);
nand gate_1389(G792,G790,G791);
nand gate_1390(G805,G803,G804);
nand gate_1391(G827,G825,G826);
nand gate_1392(G853,G851,G852);
nand gate_1393(G895,G893,G894);
nand gate_1394(G1026,G1024,G1025);
nand gate_1395(G1038,G1036,G1037);
nand gate_1396(G1055,G1053,G1054);
nand gate_1397(G1074,G1072,G1073);
nand gate_1398(G1093,G1091,G1092);
not gate_1399(G1155,G1154);
nand gate_1400(G1217,G1215,G1216);
nand gate_1401(G1226,G1224,G1225);
nand gate_1402(G1235,G1233,G1234);
nand gate_1403(G1240,G1238,G1239);
nand gate_1404(G1249,G1247,G1248);
nand gate_1405(G1258,G1256,G1257);
nand gate_1406(G1263,G1261,G1262);
nand gate_1407(G1272,G1270,G1271);
nand gate_1408(G1281,G1279,G1280);
not gate_1409(G5376,G5372);
not gate_1410(G5384,G5380);
nand gate_1411(G1546,G1544,G1545);
nand gate_1412(G1556,G1554,G1555);
nand gate_1413(G1573,G1571,G1572);
nand gate_1414(G1598,G1596,G1597);
nand gate_1415(G1609,G1607,G1608);
nand gate_1416(G1630,G1628,G1629);
nand gate_1417(G1655,G1653,G1654);
nand gate_1418(G1687,G1685,G1686);
nand gate_1419(G1695,G1693,G1694);
nand gate_1420(G1795,G1793,G1794);
nand gate_1421(G1805,G1803,G1804);
nand gate_1422(G1822,G1820,G1821);
nand gate_1423(G1850,G1848,G1849);
nand gate_1424(G1859,G1857,G1858);
nand gate_1425(G1869,G1867,G1868);
nand gate_1426(G1885,G1883,G1884);
nand gate_1427(G1903,G1901,G1902);
nand gate_1428(G1921,G1919,G1920);
not gate_1429(G5863,G5857);
nand gate_1430(G2341,G5868,G5871);
not gate_1431(G5872,G5868);
nand gate_1432(G2352,G5876,G5879);
not gate_1433(G5880,G5876);
nand gate_1434(G2370,G5884,G5887);
not gate_1435(G5888,G5884);
nand gate_1436(G2398,G5892,G5895);
not gate_1437(G5896,G5892);
nand gate_1438(G2407,G5900,G5903);
not gate_1439(G5904,G5900);
nand gate_1440(G2418,G5908,G5911);
not gate_1441(G5912,G5908);
nand gate_1442(G2434,G5916,G5919);
not gate_1443(G5920,G5916);
nand gate_1444(G2452,G5924,G5927);
not gate_1445(G5928,G5924);
and gate_1446(G2481,G3682,G4389);
not gate_1447(G5975,G5969);
nand gate_1448(G2587,G5988,G5991);
not gate_1449(G5992,G5988);
nand gate_1450(G2598,G5996,G5999);
not gate_1451(G6000,G5996);
nand gate_1452(G2616,G6004,G6007);
not gate_1453(G6008,G6004);
nand gate_1454(G2641,G6012,G6015);
not gate_1455(G6016,G6012);
nand gate_1456(G2653,G6020,G6023);
not gate_1457(G6024,G6020);
nand gate_1458(G2674,G6028,G6031);
not gate_1459(G6032,G6028);
nand gate_1460(G2699,G6036,G6039);
not gate_1461(G6040,G6036);
and gate_1462(G2724,G3682,G4389);
nand gate_1463(G2732,G6044,G6047);
not gate_1464(G6048,G6044);
nand gate_1465(G2956,G2954,G2955);
nand gate_1466(G2965,G2963,G2964);
nand gate_1467(G2973,G2971,G2972);
nand gate_1468(G2982,G2980,G2981);
nand gate_1469(G2992,G2990,G2991);
nand gate_1470(G3001,G2999,G3000);
nand gate_1471(G3009,G3007,G3008);
nand gate_1472(G3018,G3016,G3017);
nand gate_1473(G3021,G3019,G3020);
not gate_1474(G6445,G6439);
nand gate_1475(G3051,G6439,G6446);
not gate_1476(G6453,G6447);
nand gate_1477(G3061,G6447,G6454);
not gate_1478(G6461,G6455);
nand gate_1479(G3070,G6455,G6462);
not gate_1480(G6469,G6463);
nand gate_1481(G3081,G6463,G6470);
not gate_1482(G6477,G6471);
not gate_1483(G6478,G6474);
not gate_1484(G6485,G6479);
not gate_1485(G6486,G6482);
not gate_1486(G6493,G6487);
not gate_1487(G6494,G6490);
not gate_1488(G6501,G6495);
nand gate_1489(G3118,G6495,G6502);
not gate_1490(G6509,G6503);
not gate_1491(G6510,G6506);
nand gate_1492(G3176,G3174,G3175);
nand gate_1493(G3186,G3184,G3185);
nand gate_1494(G3195,G3193,G3194);
nand gate_1495(G3203,G3201,G3202);
nand gate_1496(G3215,G3213,G3214);
nand gate_1497(G3281,G6570,G6573);
not gate_1498(G6574,G6570);
nand gate_1499(G3293,G6578,G6581);
not gate_1500(G6582,G6578);
nand gate_1501(G3312,G6586,G6589);
not gate_1502(G6590,G6586);
nand gate_1503(G3342,G6594,G6597);
not gate_1504(G6598,G6594);
nand gate_1505(G3351,G6602,G6605);
not gate_1506(G6606,G6602);
nand gate_1507(G3363,G6610,G6613);
not gate_1508(G6614,G6610);
nand gate_1509(G3379,G6618,G6621);
not gate_1510(G6622,G6618);
nand gate_1511(G3397,G6626,G6629);
not gate_1512(G6630,G6626);
nand gate_1513(G3415,G6634,G6637);
not gate_1514(G6638,G6634);
not gate_1515(G6677,G6671);
nand gate_1516(G3504,G3502,G3503);
nand gate_1517(G3513,G3511,G3512);
nand gate_1518(G3522,G3520,G3521);
not gate_1519(G6727,G6721);
nand gate_1520(G3526,G6721,G6728);
not gate_1521(G6735,G6729);
not gate_1522(G6736,G6732);
not gate_1523(G6743,G6737);
not gate_1524(G6744,G6740);
not gate_1525(G6771,G6765);
nand gate_1526(G3549,G6765,G6772);
not gate_1527(G6779,G6773);
not gate_1528(G6780,G6776);
not gate_1529(G6787,G6781);
not gate_1530(G6788,G6784);
not gate_1531(G6836,G6832);
nand gate_1532(G3843,G6856,G6859);
not gate_1533(G6860,G6856);
nand gate_1534(G3854,G6864,G6867);
not gate_1535(G6868,G6864);
nand gate_1536(G3872,G6872,G6875);
not gate_1537(G6876,G6872);
nand gate_1538(G3897,G6880,G6883);
not gate_1539(G6884,G6880);
nand gate_1540(G3909,G6888,G6891);
not gate_1541(G6892,G6888);
nand gate_1542(G3930,G6896,G6899);
not gate_1543(G6900,G6896);
nand gate_1544(G3955,G6904,G6907);
not gate_1545(G6908,G6904);
nand gate_1546(G3987,G6912,G6915);
not gate_1547(G6916,G6912);
nand gate_1548(G3995,G6920,G6923);
not gate_1549(G6924,G6920);
not gate_1550(G7211,G7205);
nand gate_1551(G4179,G7205,G7212);
not gate_1552(G7219,G7213);
not gate_1553(G7220,G7216);
nand gate_1554(G4196,G7224,G7227);
not gate_1555(G7228,G7224);
nand gate_1556(G4203,G4201,G4202);
nand gate_1557(G4212,G4210,G4211);
not gate_1558(G7271,G7265);
nand gate_1559(G4220,G7265,G7272);
nand gate_1560(G4226,G4224,G4225);
nand gate_1561(G4235,G4233,G4234);
nand gate_1562(G4244,G4242,G4243);
not gate_1563(G7367,G7361);
not gate_1564(G7368,G7364);
not gate_1565(G7375,G7369);
not gate_1566(G7376,G7372);
not gate_1567(G7383,G7377);
not gate_1568(G7384,G7380);
not gate_1569(G7391,G7385);
not gate_1570(G7392,G7388);
not gate_1571(G7399,G7393);
nand gate_1572(G4326,G7393,G7400);
not gate_1573(G7407,G7401);
nand gate_1574(G4335,G7401,G7408);
not gate_1575(G7415,G7409);
nand gate_1576(G4343,G7409,G7416);
not gate_1577(G7423,G7417);
not gate_1578(G7424,G7420);
nand gate_1579(G4353,G7428,G7431);
not gate_1580(G7432,G7428);
nand gate_1581(G4531,G4529,G4530);
nand gate_1582(G4540,G4538,G4539);
nand gate_1583(G4549,G4547,G4548);
nand gate_1584(G4554,G4552,G4553);
not gate_1585(G7521,G7515);
not gate_1586(G7522,G7518);
not gate_1587(G7529,G7523);
not gate_1588(G7530,G7526);
not gate_1589(G7557,G7551);
nand gate_1590(G4576,G7551,G7558);
not gate_1591(G7565,G7559);
not gate_1592(G7566,G7562);
not gate_1593(G7573,G7567);
not gate_1594(G7574,G7570);
not gate_1595(G4936,G4932);
nand gate_1596(G4937,G4932,G4935);
not gate_1597(G4977,G4973);
nand gate_1598(G4978,G4973,G4976);
not gate_1599(G5105,G5099);
nand gate_1600(G5359,G5357,G5358);
nand gate_1601(G5362,G5347,G5348);
not gate_1602(G5529,G5523);
not gate_1603(G5675,G5669);
buf gate_1604(G5932,G4389);
buf gate_1605(G5977,G2391);
buf gate_1606(G6052,G4389);
not gate_1607(G6063,G6057);
buf gate_1608(G6115,G2635);
nor gate_1609(G6173,G3682,G4389);
buf gate_1610(G6679,G3335);
not gate_1611(G6751,G6745);
not gate_1612(G6752,G6748);
not gate_1613(G6761,G6755);
not gate_1614(G6762,G6758);
not gate_1615(G6795,G6789);
not gate_1616(G6796,G6792);
not gate_1617(G6805,G6799);
not gate_1618(G6806,G6802);
not gate_1619(G6931,G6925);
buf gate_1620(G6983,G3891);
not gate_1621(G7047,G7041);
buf gate_1622(G7129,G3979);
not gate_1623(G7279,G7273);
not gate_1624(G7280,G7276);
not gate_1625(G7289,G7283);
not gate_1626(G7290,G7286);
nand gate_1627(G7337,G7247,G7248);
nand gate_1628(G7340,G7237,G7238);
nand gate_1629(G7353,G7335,G7336);
nand gate_1630(G7356,G7325,G7326);
not gate_1631(G7537,G7531);
not gate_1632(G7538,G7534);
not gate_1633(G7547,G7541);
not gate_1634(G7548,G7544);
not gate_1635(G7581,G7575);
not gate_1636(G7582,G7578);
not gate_1637(G7591,G7585);
not gate_1638(G7592,G7588);
nand gate_1639(G7595,G7505,G7506);
nand gate_1640(G7598,G7495,G7496);
nand gate_1641(G2342,G5865,G5872);
nand gate_1642(G2353,G5873,G5880);
nand gate_1643(G2371,G5881,G5888);
nand gate_1644(G2399,G5889,G5896);
nand gate_1645(G2408,G5897,G5904);
nand gate_1646(G2419,G5905,G5912);
nand gate_1647(G2435,G5913,G5920);
nand gate_1648(G2453,G5921,G5928);
nand gate_1649(G2588,G5985,G5992);
nand gate_1650(G2599,G5993,G6000);
nand gate_1651(G2617,G6001,G6008);
nand gate_1652(G2642,G6009,G6016);
nand gate_1653(G2654,G6017,G6024);
nand gate_1654(G2675,G6025,G6032);
nand gate_1655(G2700,G6033,G6040);
nand gate_1656(G2733,G6041,G6048);
nand gate_1657(G3050,G6442,G6445);
nand gate_1658(G3060,G6450,G6453);
nand gate_1659(G3069,G6458,G6461);
nand gate_1660(G3080,G6466,G6469);
nand gate_1661(G3091,G6474,G6477);
nand gate_1662(G3092,G6471,G6478);
nand gate_1663(G3100,G6482,G6485);
nand gate_1664(G3101,G6479,G6486);
nand gate_1665(G3108,G6490,G6493);
nand gate_1666(G3109,G6487,G6494);
nand gate_1667(G3117,G6498,G6501);
nand gate_1668(G3120,G6506,G6509);
nand gate_1669(G3121,G6503,G6510);
nand gate_1670(G3282,G6567,G6574);
nand gate_1671(G3294,G6575,G6582);
nand gate_1672(G3313,G6583,G6590);
nand gate_1673(G3343,G6591,G6598);
nand gate_1674(G3352,G6599,G6606);
nand gate_1675(G3364,G6607,G6614);
nand gate_1676(G3380,G6615,G6622);
nand gate_1677(G3398,G6623,G6630);
nand gate_1678(G3416,G6631,G6638);
nand gate_1679(G3525,G6724,G6727);
nand gate_1680(G3534,G6732,G6735);
nand gate_1681(G3535,G6729,G6736);
nand gate_1682(G3543,G6740,G6743);
nand gate_1683(G3544,G6737,G6744);
nand gate_1684(G3548,G6768,G6771);
nand gate_1685(G3557,G6776,G6779);
nand gate_1686(G3558,G6773,G6780);
nand gate_1687(G3566,G6784,G6787);
nand gate_1688(G3567,G6781,G6788);
nand gate_1689(G3844,G6853,G6860);
nand gate_1690(G3855,G6861,G6868);
nand gate_1691(G3873,G6869,G6876);
nand gate_1692(G3898,G6877,G6884);
nand gate_1693(G3910,G6885,G6892);
nand gate_1694(G3931,G6893,G6900);
nand gate_1695(G3956,G6901,G6908);
nand gate_1696(G3988,G6909,G6916);
nand gate_1697(G3996,G6917,G6924);
nand gate_1698(G4178,G7208,G7211);
nand gate_1699(G4187,G7216,G7219);
nand gate_1700(G4188,G7213,G7220);
nand gate_1701(G4197,G7221,G7228);
nand gate_1702(G4219,G7268,G7271);
nand gate_1703(G4289,G7364,G7367);
nand gate_1704(G4290,G7361,G7368);
nand gate_1705(G4298,G7372,G7375);
nand gate_1706(G4299,G7369,G7376);
nand gate_1707(G4306,G7380,G7383);
nand gate_1708(G4307,G7377,G7384);
nand gate_1709(G4315,G7388,G7391);
nand gate_1710(G4316,G7385,G7392);
nand gate_1711(G4325,G7396,G7399);
nand gate_1712(G4334,G7404,G7407);
nand gate_1713(G4342,G7412,G7415);
nand gate_1714(G4350,G7420,G7423);
nand gate_1715(G4351,G7417,G7424);
nand gate_1716(G4354,G7425,G7432);
nand gate_1717(G4561,G7518,G7521);
nand gate_1718(G4562,G7515,G7522);
nand gate_1719(G4570,G7526,G7529);
nand gate_1720(G4571,G7523,G7530);
nand gate_1721(G4575,G7554,G7557);
nand gate_1722(G4584,G7562,G7565);
nand gate_1723(G4585,G7559,G7566);
nand gate_1724(G4593,G7570,G7573);
nand gate_1725(G4594,G7567,G7574);
nand gate_1726(G4938,G4929,G4936);
nand gate_1727(G4979,G4970,G4977);
nand gate_1728(G6753,G6748,G6751);
nand gate_1729(G6754,G6745,G6752);
nand gate_1730(G6763,G6758,G6761);
nand gate_1731(G6764,G6755,G6762);
nand gate_1732(G6797,G6792,G6795);
nand gate_1733(G6798,G6789,G6796);
nand gate_1734(G6807,G6802,G6805);
nand gate_1735(G6808,G6799,G6806);
nand gate_1736(G7281,G7276,G7279);
nand gate_1737(G7282,G7273,G7280);
nand gate_1738(G7291,G7286,G7289);
nand gate_1739(G7292,G7283,G7290);
nand gate_1740(G7539,G7534,G7537);
nand gate_1741(G7540,G7531,G7538);
nand gate_1742(G7549,G7544,G7547);
nand gate_1743(G7550,G7541,G7548);
nand gate_1744(G7583,G7578,G7581);
nand gate_1745(G7584,G7575,G7582);
nand gate_1746(G7593,G7588,G7591);
nand gate_1747(G7594,G7585,G7592);
not gate_1748(G1856,G1850);
and gate_1749(G920,G895,G853,G827,G805,G792);
and gate_1750(G925,G792,G821);
and gate_1751(G926,G805,G792,G845);
and gate_1752(G927,G827,G792,G868,G805);
and gate_1753(G928,G853,G827,G792,G877,G805);
and gate_1754(G937,G805,G845);
and gate_1755(G938,G827,G868,G805);
and gate_1756(G939,G853,G827,G877,G805);
and gate_1757(G940,G895,G827,G805,G853);
and gate_1758(G941,G805,G845);
and gate_1759(G942,G827,G868,G805);
and gate_1760(G943,G853,G827,G877,G805);
and gate_1761(G944,G827,G868);
and gate_1762(G945,G853,G827,G877);
and gate_1763(G946,G895,G827,G853);
and gate_1764(G947,G827,G868);
and gate_1765(G948,G853,G827,G877);
and gate_1766(G949,G853,G877);
and gate_1767(G956,G895,G853);
and gate_1768(G1122,G1038,G1093,G1055,G1026,G1074);
and gate_1769(G1125,G1026,G1050);
and gate_1770(G1126,G1038,G1026,G1068);
and gate_1771(G1127,G1055,G1026,G1086,G1038);
and gate_1772(G1128,G1074,G1055,G1026,G1102,G1038);
and gate_1773(G1132,G1038,G1068);
and gate_1774(G1133,G1055,G1086,G1038);
and gate_1775(G1134,G1074,G1055,G1102,G1038);
and gate_1776(G1137,G1086,G1055);
and gate_1777(G1138,G1074,G1055,G1102);
and gate_1778(G1141,G1074,G1102);
not gate_1779(G1221,G1217);
not gate_1780(G1230,G1226);
not gate_1781(G1244,G1240);
not gate_1782(G1253,G1249);
not gate_1783(G1267,G1263);
not gate_1784(G1276,G1272);
buf gate_1785(G1284,G1235);
buf gate_1786(G1288,G1235);
buf gate_1787(G1292,G1258);
buf gate_1788(G1296,G1258);
buf gate_1789(G1300,G1281);
buf gate_1790(G1304,G1281);
and gate_1791(G1702,G1687,G1573,G1556,G1546);
and gate_1792(G1705,G1546,G1567);
and gate_1793(G1706,G1556,G1546,G1584);
and gate_1794(G1707,G1573,G1546,G1590,G1556);
and gate_1795(G1709,G1556,G1584);
and gate_1796(G1710,G1573,G1590,G1556);
and gate_1797(G1711,G1687,G1573,G1556);
and gate_1798(G1712,G1556,G1584);
and gate_1799(G1713,G1573,G1590,G1556);
and gate_1800(G1714,G1573,G1590);
and gate_1801(G1718,G1695,G1655,G1630,G1609,G1598);
and gate_1802(G1722,G1598,G1624);
and gate_1803(G1723,G1609,G1598,G1647);
and gate_1804(G1724,G1630,G1598,G1669,G1609);
and gate_1805(G1725,G1655,G1630,G1598,G1677,G1609);
and gate_1806(G1733,G1609,G1647);
and gate_1807(G1734,G1630,G1669,G1609);
and gate_1808(G1735,G1655,G1630,G1677,G1609);
and gate_1809(G1736,G1695,G1630,G1609,G1655);
and gate_1810(G1737,G1609,G1647);
and gate_1811(G1738,G1630,G1669,G1609);
and gate_1812(G1739,G1655,G1630,G1677,G1609);
and gate_1813(G1740,G1630,G1669);
and gate_1814(G1741,G1655,G1630,G1677);
and gate_1815(G1742,G1695,G1630,G1655);
and gate_1816(G1743,G1630,G1669);
and gate_1817(G1744,G1655,G1630,G1677);
and gate_1818(G1745,G1655,G1677);
and gate_1819(G1749,G1687,G1573);
and gate_1820(G1750,G1695,G1655);
and gate_1821(G1935,G1805,G1850,G1822,G1795);
and gate_1822(G1938,G1795,G1816);
and gate_1823(G1939,G1805,G1795,G1834);
and gate_1824(G1940,G1822,G1795,G1841,G1805);
and gate_1825(G1942,G1805,G1834);
and gate_1826(G1943,G1822,G1841,G1805);
and gate_1827(G1944,G1850,G1822,G1805);
and gate_1828(G1945,G1805,G1834);
and gate_1829(G1946,G1841,G1822,G1805);
and gate_1830(G1947,G1822,G1841);
and gate_1831(G1948,G1850,G1822);
and gate_1832(G1949,G1822,G1841);
and gate_1833(G1950,G1869,G1921,G1885,G1859,G1903);
and gate_1834(G1953,G1859,G1880);
and gate_1835(G1954,G1869,G1859,G1897);
and gate_1836(G1955,G1885,G1859,G1914,G1869);
and gate_1837(G1956,G1903,G1885,G1859,G1929,G1869);
and gate_1838(G1960,G1869,G1897);
and gate_1839(G1961,G1885,G1914,G1869);
and gate_1840(G1962,G1903,G1885,G1929,G1869);
and gate_1841(G1965,G1914,G1885);
and gate_1842(G1966,G1903,G1885,G1929);
and gate_1843(G1969,G1903,G1929);
nand gate_1844(G2343,G2341,G2342);
nand gate_1845(G2354,G2352,G2353);
nand gate_1846(G2372,G2370,G2371);
nand gate_1847(G2400,G2398,G2399);
nand gate_1848(G2409,G2407,G2408);
nand gate_1849(G2420,G2418,G2419);
nand gate_1850(G2436,G2434,G2435);
nand gate_1851(G2454,G2452,G2453);
nand gate_1852(G2470,G5932,G5935);
not gate_1853(G5936,G5932);
not gate_1854(G5983,G5977);
nand gate_1855(G2589,G2587,G2588);
nand gate_1856(G2600,G2598,G2599);
nand gate_1857(G2618,G2616,G2617);
nand gate_1858(G2643,G2641,G2642);
nand gate_1859(G2655,G2653,G2654);
nand gate_1860(G2676,G2674,G2675);
nand gate_1861(G2701,G2699,G2700);
nand gate_1862(G2734,G2732,G2733);
nand gate_1863(G2740,G6052,G6055);
not gate_1864(G6056,G6052);
and gate_1865(G3022,G3018,G2973,G2965,G2956);
and gate_1866(G3025,G2956,G2970);
and gate_1867(G3026,G2965,G2956,G2977);
and gate_1868(G3027,G2973,G2956,G2979,G2965);
and gate_1869(G3029,G3021,G3009,G3001,G2992,G2982);
and gate_1870(G3030,G2982,G2998);
and gate_1871(G3031,G2992,G2982,G3006);
and gate_1872(G3032,G3001,G2982,G3013,G2992);
and gate_1873(G3033,G3009,G3001,G2982,G3015,G2992);
nand gate_1874(G3052,G3050,G3051);
nand gate_1875(G3062,G3060,G3061);
nand gate_1876(G3071,G3069,G3070);
nand gate_1877(G3082,G3080,G3081);
nand gate_1878(G3093,G3091,G3092);
nand gate_1879(G3102,G3100,G3101);
nand gate_1880(G3110,G3108,G3109);
nand gate_1881(G3119,G3117,G3118);
nand gate_1882(G3122,G3120,G3121);
and gate_1883(G3228,G3215,G3203,G3195,G3186,G3176);
and gate_1884(G3231,G3176,G3192);
and gate_1885(G3232,G3186,G3176,G3200);
and gate_1886(G3233,G3195,G3176,G3207,G3186);
and gate_1887(G3234,G3203,G3195,G3176,G3209,G3186);
nand gate_1888(G3283,G3281,G3282);
nand gate_1889(G3295,G3293,G3294);
nand gate_1890(G3314,G3312,G3313);
nand gate_1891(G3344,G3342,G3343);
nand gate_1892(G3353,G3351,G3352);
nand gate_1893(G3365,G3363,G3364);
nand gate_1894(G3381,G3379,G3380);
nand gate_1895(G3399,G3397,G3398);
nand gate_1896(G3417,G3415,G3416);
not gate_1897(G6685,G6679);
not gate_1898(G3508,G3504);
not gate_1899(G3517,G3513);
nand gate_1900(G3527,G3525,G3526);
nand gate_1901(G3536,G3534,G3535);
nand gate_1902(G3545,G3543,G3544);
nand gate_1903(G3550,G3548,G3549);
nand gate_1904(G3559,G3557,G3558);
nand gate_1905(G3568,G3566,G3567);
buf gate_1906(G3571,G3522);
buf gate_1907(G3575,G3522);
nand gate_1908(G3845,G3843,G3844);
nand gate_1909(G3856,G3854,G3855);
nand gate_1910(G3874,G3872,G3873);
nand gate_1911(G3899,G3897,G3898);
nand gate_1912(G3911,G3909,G3910);
nand gate_1913(G3932,G3930,G3931);
nand gate_1914(G3957,G3955,G3956);
nand gate_1915(G3989,G3987,G3988);
nand gate_1916(G3997,G3995,G3996);
nand gate_1917(G4180,G4178,G4179);
nand gate_1918(G4189,G4187,G4188);
nand gate_1919(G4198,G4196,G4197);
not gate_1920(G4207,G4203);
not gate_1921(G4216,G4212);
nand gate_1922(G4221,G4219,G4220);
not gate_1923(G4230,G4226);
not gate_1924(G4239,G4235);
buf gate_1925(G4263,G4244);
buf gate_1926(G4267,G4244);
nand gate_1927(G4291,G4289,G4290);
nand gate_1928(G4300,G4298,G4299);
nand gate_1929(G4308,G4306,G4307);
nand gate_1930(G4317,G4315,G4316);
nand gate_1931(G4327,G4325,G4326);
nand gate_1932(G4336,G4334,G4335);
nand gate_1933(G4344,G4342,G4343);
nand gate_1934(G4352,G4350,G4351);
nand gate_1935(G4355,G4353,G4354);
not gate_1936(G4535,G4531);
not gate_1937(G4544,G4540);
not gate_1938(G4558,G4554);
nand gate_1939(G4563,G4561,G4562);
nand gate_1940(G4572,G4570,G4571);
nand gate_1941(G4577,G4575,G4576);
nand gate_1942(G4586,G4584,G4585);
nand gate_1943(G4595,G4593,G4594);
buf gate_1944(G4598,G4549);
buf gate_1945(G4602,G4549);
buf gate_1946(G4716,G1921);
buf gate_1947(G4724,G1859);
buf gate_1948(G4732,G1869);
buf gate_1949(G4740,G1885);
buf gate_1950(G4748,G1903);
buf gate_1951(G4756,G1093);
buf gate_1952(G4764,G1026);
buf gate_1953(G4772,G1038);
buf gate_1954(G4780,G1055);
buf gate_1955(G4788,G1074);
nand gate_1956(G4939,G4937,G4938);
nand gate_1957(G4980,G4978,G4979);
buf gate_1958(G5044,G895);
buf gate_1959(G5054,G853);
buf gate_1960(G5064,G792);
buf gate_1961(G5074,G827);
buf gate_1962(G5084,G805);
buf gate_1963(G5094,G805);
buf gate_1964(G5132,G895);
buf gate_1965(G5142,G853);
buf gate_1966(G5152,G792);
buf gate_1967(G5162,G827);
not gate_1968(G5365,G5359);
not gate_1969(G5366,G5362);
buf gate_1970(G5488,G1687);
buf gate_1971(G5498,G1573);
buf gate_1972(G5508,G1546);
buf gate_1973(G5518,G1556);
buf gate_1974(G5546,G1687);
buf gate_1975(G5556,G1573);
buf gate_1976(G5566,G1546);
buf gate_1977(G5576,G1556);
buf gate_1978(G5614,G1695);
buf gate_1979(G5624,G1655);
buf gate_1980(G5634,G1598);
buf gate_1981(G5644,G1630);
buf gate_1982(G5654,G1609);
buf gate_1983(G5664,G1609);
buf gate_1984(G5702,G1695);
buf gate_1985(G5712,G1655);
buf gate_1986(G5722,G1598);
buf gate_1987(G5732,G1630);
buf gate_1988(G5820,G1795);
buf gate_1989(G5828,G1795);
buf gate_1990(G5836,G1805);
buf gate_1991(G5844,G1805);
buf gate_1992(G5852,G1822);
buf gate_1993(G5860,G1822);
not gate_1994(G6121,G6115);
not gate_1995(G6179,G6173);
buf gate_1996(G6261,G2724);
not gate_1997(G7359,G7353);
not gate_1998(G7360,G7356);
not gate_1999(G7343,G7337);
not gate_2000(G7344,G7340);
nand gate_2001(G6809,G6763,G6764);
nand gate_2002(G6812,G6753,G6754);
nand gate_2003(G6819,G6807,G6808);
nand gate_2004(G6822,G6797,G6798);
not gate_2005(G6989,G6983);
not gate_2006(G7135,G7129);
nand gate_2007(G7345,G7291,G7292);
nand gate_2008(G7348,G7281,G7282);
not gate_2009(G7601,G7595);
not gate_2010(G7602,G7598);
nand gate_2011(G7603,G7549,G7550);
nand gate_2012(G7606,G7539,G7540);
nand gate_2013(G7611,G7593,G7594);
nand gate_2014(G7614,G7583,G7584);
or gate_2015(G929,G802,G925,G926,G927,G928);
or gate_2016(G950,G868,G949);
or gate_2017(G1129,G1035,G1125,G1126,G1127,G1128);
or gate_2018(G1708,G1553,G1705,G1706,G1707);
or gate_2019(G1715,G1584,G1714);
or gate_2020(G1726,G1606,G1722,G1723,G1724,G1725);
or gate_2021(G1746,G1669,G1745);
or gate_2022(G1941,G1802,G1938,G1939,G1940);
or gate_2023(G1957,G1866,G1953,G1954,G1955,G1956);
nand gate_2024(G2471,G5929,G5936);
nand gate_2025(G2741,G6049,G6056);
or gate_2026(G3028,G2962,G3025,G3026,G3027);
or gate_2027(G3034,G2989,G3030,G3031,G3032,G3033);
or gate_2028(G3235,G3183,G3231,G3232,G3233,G3234);
or gate_2029(G5014,G845,G944,G945,G946);
or gate_2030(G5034,G821,G937,G938,G939,G940);
nor gate_2031(G5102,G845,G947,G948);
nor gate_2032(G5122,G821,G941,G942,G943);
nand gate_2033(G5367,G5362,G5365);
nand gate_2034(G5368,G5359,G5366);
or gate_2035(G5478,G1567,G1709,G1710,G1711);
nor gate_2036(G5536,G1567,G1712,G1713);
or gate_2037(G5584,G1647,G1740,G1741,G1742);
or gate_2038(G5604,G1624,G1733,G1734,G1735,G1736);
nor gate_2039(G5672,G1647,G1743,G1744);
nor gate_2040(G5692,G1624,G1737,G1738,G1739);
or gate_2041(G5817,G1816,G1942,G1943,G1944);
nor gate_2042(G5825,G1816,G1945,G1946);
or gate_2043(G5833,G1834,G1947,G1948);
nor gate_2044(G5841,G1834,G1949);
nand gate_2045(G6340,G7356,G7359);
nand gate_2046(G6341,G7353,G7360);
nand gate_2047(G6350,G7340,G7343);
nand gate_2048(G6351,G7337,G7344);
nand gate_2049(G7436,G7598,G7601);
nand gate_2050(G7437,G7595,G7602);
not gate_2051(G4720,G4716);
not gate_2052(G4728,G4724);
not gate_2053(G4736,G4732);
not gate_2054(G4744,G4740);
not gate_2055(G4752,G4748);
not gate_2056(G4760,G4756);
not gate_2057(G4768,G4764);
not gate_2058(G4776,G4772);
not gate_2059(G4784,G4780);
not gate_2060(G4792,G4788);
not gate_2061(G3350,G3344);
not gate_2062(G2406,G2400);
not gate_2063(G924,G920);
not gate_2064(G5088,G5084);
not gate_2065(G5098,G5094);
and gate_2066(G997,G902,G920);
and gate_2067(G1146,G1108,G1122);
not gate_2068(G1287,G1284);
not gate_2069(G1291,G1288);
not gate_2070(G1295,G1292);
not gate_2071(G1299,G1296);
not gate_2072(G1303,G1300);
not gate_2073(G1307,G1304);
and gate_2074(G1309,G1226,G1217,G1284);
and gate_2075(G1312,G1230,G1221,G1288);
and gate_2076(G1315,G1249,G1240,G1292);
and gate_2077(G1318,G1253,G1244,G1296);
and gate_2078(G1321,G1272,G1263,G1300);
and gate_2079(G1324,G1276,G1267,G1304);
not gate_2080(G1721,G1718);
not gate_2081(G5522,G5518);
not gate_2082(G5580,G5576);
not gate_2083(G5658,G5654);
not gate_2084(G5668,G5664);
and gate_2085(G1788,G1702,G1718);
and gate_2086(G1974,G1935,G1950);
not gate_2087(G5824,G5820);
not gate_2088(G5832,G5828);
not gate_2089(G5840,G5836);
not gate_2090(G5848,G5844);
nand gate_2091(G1999,G5852,G5855);
not gate_2092(G5856,G5852);
nand gate_2093(G2003,G5860,G5863);
not gate_2094(G5864,G5860);
nand gate_2095(G2472,G2470,G2471);
and gate_2096(G2487,G2354,G2400,G2372,G2343);
and gate_2097(G2492,G2343,G2366);
and gate_2098(G2493,G2354,G2343,G2384);
and gate_2099(G2494,G2372,G2343,G2391,G2354);
and gate_2100(G2500,G2354,G2384);
and gate_2101(G2501,G2372,G2391,G2354);
and gate_2102(G2502,G2400,G2372,G2354);
and gate_2103(G2503,G2354,G2384);
and gate_2104(G2504,G2391,G2372,G2354);
and gate_2105(G2505,G2372,G2391);
and gate_2106(G2506,G2400,G2372);
and gate_2107(G2507,G2372,G2391);
and gate_2108(G2511,G2409,G2431);
and gate_2109(G2512,G2420,G2409,G2448);
and gate_2110(G2513,G2436,G2409,G2465,G2420);
and gate_2111(G2514,G2454,G2436,G2409,G2481,G2420);
and gate_2112(G2518,G2420,G2448);
and gate_2113(G2519,G2436,G2465,G2420);
and gate_2114(G2520,G2454,G2436,G2481,G2420);
and gate_2115(G2523,G2465,G2436);
and gate_2116(G2524,G2454,G2436,G2481);
and gate_2117(G2527,G2454,G2481);
nand gate_2118(G2742,G2740,G2741);
and gate_2119(G2749,G2734,G2618,G2600,G2589);
and gate_2120(G2754,G2589,G2612);
and gate_2121(G2755,G2600,G2589,G2629);
and gate_2122(G2756,G2618,G2589,G2635,G2600);
and gate_2123(G2762,G2600,G2629);
and gate_2124(G2763,G2618,G2635,G2600);
and gate_2125(G2764,G2734,G2618,G2600);
and gate_2126(G2765,G2600,G2629);
and gate_2127(G2766,G2618,G2635,G2600);
and gate_2128(G2767,G2618,G2635);
and gate_2129(G2776,G2643,G2670);
and gate_2130(G2777,G2655,G2643,G2693);
and gate_2131(G2778,G2676,G2643,G2715,G2655);
and gate_2132(G2779,G2701,G2676,G2643,G2724,G2655);
and gate_2133(G2788,G2655,G2693);
and gate_2134(G2789,G2676,G2715,G2655);
and gate_2135(G2790,G2701,G2676,G2724,G2655);
and gate_2136(G2792,G2655,G2693);
and gate_2137(G2793,G2676,G2715,G2655);
and gate_2138(G2794,G2701,G2676,G2724,G2655);
and gate_2139(G2795,G2676,G2715);
and gate_2140(G2796,G2701,G2676,G2724);
and gate_2141(G2798,G2676,G2715);
and gate_2142(G2799,G2701,G2676,G2724);
and gate_2143(G2800,G2701,G2724);
and gate_2144(G2804,G2734,G2618);
and gate_2145(G3035,G3022,G3029);
and gate_2146(G3045,G3022,G3034);
and gate_2147(G3123,G3119,G3071,G3062,G3052);
and gate_2148(G3128,G3052,G3068);
and gate_2149(G3129,G3062,G3052,G3076);
and gate_2150(G3130,G3071,G3052,G3079,G3062);
and gate_2151(G3136,G3122,G3110,G3102,G3093,G3082);
and gate_2152(G3139,G3082,G3099);
and gate_2153(G3140,G3093,G3082,G3107);
and gate_2154(G3141,G3102,G3082,G3114,G3093);
and gate_2155(G3142,G3110,G3102,G3082,G3116,G3093);
and gate_2156(G3249,G3216,G3228);
and gate_2157(G3431,G3295,G3344,G3314,G3283);
and gate_2158(G3434,G3283,G3308);
and gate_2159(G3435,G3295,G3283,G3327);
and gate_2160(G3436,G3314,G3283,G3335,G3295);
and gate_2161(G3438,G3295,G3327);
and gate_2162(G3439,G3314,G3335,G3295);
and gate_2163(G3440,G3344,G3314,G3295);
and gate_2164(G3441,G3295,G3327);
and gate_2165(G3442,G3335,G3314,G3295);
and gate_2166(G3443,G3314,G3335);
and gate_2167(G3444,G3344,G3314);
and gate_2168(G3445,G3314,G3335);
and gate_2169(G3446,G3365,G3417,G3381,G3353,G3399);
and gate_2170(G3449,G3353,G3376);
and gate_2171(G3450,G3365,G3353,G3393);
and gate_2172(G3451,G3381,G3353,G3410,G3365);
and gate_2173(G3452,G3399,G3381,G3353,G3425,G3365);
and gate_2174(G3456,G3365,G3393);
and gate_2175(G3457,G3381,G3410,G3365);
and gate_2176(G3458,G3399,G3381,G3425,G3365);
and gate_2177(G3460,G3410,G3381);
and gate_2178(G3461,G3399,G3381,G3425);
and gate_2179(G3463,G3399,G3425);
not gate_2180(G3531,G3527);
not gate_2181(G3540,G3536);
not gate_2182(G3554,G3550);
not gate_2183(G3563,G3559);
not gate_2184(G3574,G3571);
not gate_2185(G3578,G3575);
buf gate_2186(G3579,G3545);
buf gate_2187(G3583,G3545);
buf gate_2188(G3587,G3568);
buf gate_2189(G3591,G3568);
and gate_2190(G3596,G3513,G3504,G3571);
and gate_2191(G3599,G3517,G3508,G3575);
and gate_2192(G4004,G3989,G3874,G3856,G3845);
and gate_2193(G4007,G3845,G3868);
and gate_2194(G4008,G3856,G3845,G3885);
and gate_2195(G4009,G3874,G3845,G3891,G3856);
and gate_2196(G4011,G3856,G3885);
and gate_2197(G4012,G3874,G3891,G3856);
and gate_2198(G4013,G3989,G3874,G3856);
and gate_2199(G4014,G3856,G3885);
and gate_2200(G4015,G3874,G3891,G3856);
and gate_2201(G4016,G3874,G3891);
and gate_2202(G4020,G3997,G3957,G3932,G3911,G3899);
and gate_2203(G4024,G3899,G3926);
and gate_2204(G4025,G3911,G3899,G3949);
and gate_2205(G4026,G3932,G3899,G3971,G3911);
and gate_2206(G4027,G3957,G3932,G3899,G3979,G3911);
and gate_2207(G4035,G3911,G3949);
and gate_2208(G4036,G3932,G3971,G3911);
and gate_2209(G4037,G3957,G3932,G3979,G3911);
and gate_2210(G4038,G3997,G3932,G3911,G3957);
and gate_2211(G4039,G3911,G3949);
and gate_2212(G4040,G3932,G3971,G3911);
and gate_2213(G4041,G3957,G3932,G3979,G3911);
and gate_2214(G4042,G3932,G3971);
and gate_2215(G4043,G3957,G3932,G3979);
and gate_2216(G4044,G3997,G3932,G3957);
and gate_2217(G4045,G3932,G3971);
and gate_2218(G4046,G3957,G3932,G3979);
and gate_2219(G4047,G3957,G3979);
and gate_2220(G4051,G3989,G3874);
and gate_2221(G4052,G3997,G3957);
not gate_2222(G4184,G4180);
not gate_2223(G4193,G4189);
buf gate_2224(G4247,G4198);
buf gate_2225(G4251,G4198);
buf gate_2226(G4255,G4221);
buf gate_2227(G4259,G4221);
not gate_2228(G4266,G4263);
not gate_2229(G4270,G4267);
and gate_2230(G4284,G4235,G4226,G4263);
and gate_2231(G4287,G4239,G4230,G4267);
and gate_2232(G4356,G4352,G4308,G4300,G4291);
and gate_2233(G4361,G4291,G4305);
and gate_2234(G4362,G4300,G4291,G4312);
and gate_2235(G4363,G4308,G4291,G4314,G4300);
and gate_2236(G4369,G4355,G4344,G4336,G4327,G4317);
and gate_2237(G4372,G4317,G4333);
and gate_2238(G4373,G4327,G4317,G4341);
and gate_2239(G4374,G4336,G4317,G4348,G4327);
and gate_2240(G4375,G4344,G4336,G4317,G4349,G4327);
not gate_2241(G4567,G4563);
not gate_2242(G4581,G4577);
not gate_2243(G4590,G4586);
not gate_2244(G4601,G4598);
not gate_2245(G4605,G4602);
buf gate_2246(G4606,G4572);
buf gate_2247(G4610,G4572);
buf gate_2248(G4614,G4595);
buf gate_2249(G4618,G4595);
and gate_2250(G4623,G4540,G4531,G4598);
and gate_2251(G4626,G4544,G4535,G4602);
buf gate_2252(G4796,G3417);
buf gate_2253(G4804,G3353);
buf gate_2254(G4812,G3365);
buf gate_2255(G4820,G3381);
buf gate_2256(G4828,G3399);
buf gate_2257(G4844,G2409);
buf gate_2258(G4852,G2420);
buf gate_2259(G4860,G2436);
buf gate_2260(G4868,G2454);
not gate_2261(G4945,G4939);
nand gate_2262(G4948,G4939,G4946);
not gate_2263(G4986,G4980);
nand gate_2264(G4989,G4980,G4987);
not gate_2265(G5048,G5044);
not gate_2266(G5058,G5054);
not gate_2267(G5068,G5064);
not gate_2268(G5078,G5074);
not gate_2269(G5166,G5162);
not gate_2270(G5136,G5132);
not gate_2271(G5146,G5142);
not gate_2272(G5156,G5152);
nand gate_2273(G5388,G5367,G5368);
not gate_2274(G5492,G5488);
not gate_2275(G5502,G5498);
not gate_2276(G5512,G5508);
not gate_2277(G5550,G5546);
not gate_2278(G5560,G5556);
not gate_2279(G5570,G5566);
not gate_2280(G5618,G5614);
not gate_2281(G5628,G5624);
not gate_2282(G5638,G5634);
not gate_2283(G5648,G5644);
not gate_2284(G5736,G5732);
not gate_2285(G5706,G5702);
not gate_2286(G5716,G5712);
not gate_2287(G5726,G5722);
buf gate_2288(G5940,G2343);
buf gate_2289(G5948,G2343);
buf gate_2290(G5956,G2354);
buf gate_2291(G5964,G2354);
buf gate_2292(G5972,G2372);
buf gate_2293(G5980,G2372);
buf gate_2294(G6080,G2734);
buf gate_2295(G6090,G2618);
buf gate_2296(G6100,G2589);
buf gate_2297(G6110,G2600);
buf gate_2298(G6138,G2734);
buf gate_2299(G6148,G2618);
buf gate_2300(G6158,G2589);
buf gate_2301(G6168,G2600);
buf gate_2302(G6216,G2701);
buf gate_2303(G6226,G2643);
buf gate_2304(G6236,G2676);
buf gate_2305(G6246,G2655);
buf gate_2306(G6256,G2655);
not gate_2307(G6267,G6261);
buf gate_2308(G6304,G2701);
buf gate_2309(G6314,G2643);
buf gate_2310(G6324,G2676);
nand gate_2311(G6342,G6340,G6341);
nand gate_2312(G6352,G6350,G6351);
not gate_2313(G7351,G7345);
not gate_2314(G7352,G7348);
buf gate_2315(G6642,G3283);
buf gate_2316(G6650,G3283);
buf gate_2317(G6658,G3295);
buf gate_2318(G6666,G3295);
buf gate_2319(G6674,G3314);
buf gate_2320(G6682,G3314);
not gate_2321(G6815,G6809);
not gate_2322(G6816,G6812);
not gate_2323(G6825,G6819);
not gate_2324(G6826,G6822);
buf gate_2325(G6948,G3989);
buf gate_2326(G6958,G3874);
buf gate_2327(G6968,G3845);
buf gate_2328(G6978,G3856);
buf gate_2329(G7006,G3989);
buf gate_2330(G7016,G3874);
buf gate_2331(G7026,G3845);
buf gate_2332(G7036,G3856);
buf gate_2333(G7074,G3997);
buf gate_2334(G7084,G3957);
buf gate_2335(G7094,G3899);
buf gate_2336(G7104,G3932);
buf gate_2337(G7114,G3911);
buf gate_2338(G7124,G3911);
buf gate_2339(G7162,G3997);
buf gate_2340(G7172,G3957);
buf gate_2341(G7182,G3899);
buf gate_2342(G7192,G3932);
nand gate_2343(G7438,G7436,G7437);
not gate_2344(G7617,G7611);
not gate_2345(G7618,G7614);
not gate_2346(G7609,G7603);
not gate_2347(G7610,G7606);
and gate_2348(G1151,G1129,G1108);
and gate_2349(G1002,G902,G929);
not gate_2350(G933,G929);
and gate_2351(G1308,G1221,G1226,G1287);
and gate_2352(G1311,G1217,G1230,G1291);
and gate_2353(G1314,G1244,G1249,G1295);
and gate_2354(G1317,G1240,G1253,G1299);
and gate_2355(G1320,G1267,G1272,G1303);
and gate_2356(G1323,G1263,G1276,G1307);
not gate_2357(G1730,G1726);
and gate_2358(G1789,G1702,G1726);
and gate_2359(G1981,G1957,G1935);
not gate_2360(G5823,G5817);
nand gate_2361(G1986,G5817,G5824);
not gate_2362(G5831,G5825);
nand gate_2363(G1989,G5825,G5832);
not gate_2364(G5839,G5833);
nand gate_2365(G1993,G5833,G5840);
not gate_2366(G5847,G5841);
nand gate_2367(G1996,G5841,G5848);
nand gate_2368(G2000,G5849,G5856);
nand gate_2369(G2004,G5857,G5864);
or gate_2370(G2495,G2351,G2492,G2493,G2494);
or gate_2371(G2515,G2417,G2511,G2512,G2513,G2514);
or gate_2372(G2757,G2597,G2754,G2755,G2756);
or gate_2373(G2768,G2629,G2767);
or gate_2374(G2780,G2652,G2776,G2777,G2778,G2779);
or gate_2375(G2801,G2715,G2800);
or gate_2376(G3046,G3028,G3045);
or gate_2377(G3131,G3059,G3128,G3129,G3130);
or gate_2378(G3143,G3090,G3139,G3140,G3141,G3142);
not gate_2379(G3238,G3235);
and gate_2380(G3258,G3216,G3235);
or gate_2381(G3437,G3292,G3434,G3435,G3436);
or gate_2382(G3453,G3362,G3449,G3450,G3451,G3452);
and gate_2383(G3595,G3508,G3513,G3574);
and gate_2384(G3598,G3504,G3517,G3578);
or gate_2385(G4010,G3853,G4007,G4008,G4009);
or gate_2386(G4017,G3885,G4016);
or gate_2387(G4028,G3908,G4024,G4025,G4026,G4027);
or gate_2388(G4048,G3971,G4047);
and gate_2389(G4283,G4230,G4235,G4266);
and gate_2390(G4286,G4226,G4239,G4270);
or gate_2391(G4364,G4297,G4361,G4362,G4363);
or gate_2392(G4376,G4324,G4372,G4373,G4374,G4375);
and gate_2393(G4622,G4535,G4540,G4601);
and gate_2394(G4625,G4531,G4544,G4605);
nand gate_2395(G4947,G4942,G4945);
nand gate_2396(G4988,G4983,G4986);
not gate_2397(G5018,G5014);
nand gate_2398(G5019,G5014,G5017);
or gate_2399(G5024,G950,G956);
not gate_2400(G5038,G5034);
not gate_2401(G5106,G5102);
nand gate_2402(G5107,G5102,G5105);
not gate_2403(G5112,G950);
not gate_2404(G5126,G5122);
or gate_2405(G5468,G1715,G1749);
not gate_2406(G5482,G5478);
not gate_2407(G5526,G1715);
not gate_2408(G5540,G5536);
not gate_2409(G5588,G5584);
nand gate_2410(G5589,G5584,G5587);
or gate_2411(G5594,G1746,G1750);
not gate_2412(G5608,G5604);
not gate_2413(G5676,G5672);
nand gate_2414(G5677,G5672,G5675);
not gate_2415(G5682,G1746);
not gate_2416(G5696,G5692);
or gate_2417(G5937,G2366,G2500,G2501,G2502);
nor gate_2418(G5945,G2366,G2503,G2504);
or gate_2419(G5953,G2384,G2505,G2506);
nor gate_2420(G5961,G2384,G2507);
or gate_2421(G6070,G2612,G2762,G2763,G2764);
nor gate_2422(G6128,G2612,G2765,G2766);
nor gate_2423(G6264,G2693,G2798,G2799);
nor gate_2424(G6284,G2670,G2792,G2793,G2794);
nand gate_2425(G6360,G7348,G7351);
nand gate_2426(G6361,G7345,G7352);
or gate_2427(G6639,G3308,G3438,G3439,G3440);
nor gate_2428(G6647,G3308,G3441,G3442);
or gate_2429(G6655,G3327,G3443,G3444);
nor gate_2430(G6663,G3327,G3445);
nand gate_2431(G6817,G6812,G6815);
nand gate_2432(G6818,G6809,G6816);
nand gate_2433(G6827,G6822,G6825);
nand gate_2434(G6828,G6819,G6826);
or gate_2435(G6938,G3868,G4011,G4012,G4013);
nor gate_2436(G6996,G3868,G4014,G4015);
or gate_2437(G7044,G3949,G4042,G4043,G4044);
or gate_2438(G7064,G3926,G4035,G4036,G4037,G4038);
nor gate_2439(G7132,G3949,G4045,G4046);
nor gate_2440(G7152,G3926,G4039,G4040,G4041);
nand gate_2441(G7446,G7614,G7617);
nand gate_2442(G7447,G7611,G7618);
nand gate_2443(G7456,G7606,G7609);
nand gate_2444(G7457,G7603,G7610);
or gate_2445(G241,G1117,G1151);
or gate_2446(G265,G908,G1002);
nand gate_2447(G2005,G2003,G2004);
not gate_2448(G4800,G4796);
not gate_2449(G4808,G4804);
not gate_2450(G4816,G4812);
not gate_2451(G4824,G4820);
not gate_2452(G4832,G4828);
not gate_2453(G4848,G4844);
not gate_2454(G4856,G4852);
not gate_2455(G4864,G4860);
not gate_2456(G4872,G4868);
nor gate_2457(G1310,G1308,G1309);
nor gate_2458(G1313,G1311,G1312);
nor gate_2459(G1316,G1314,G1315);
nor gate_2460(G1319,G1317,G1318);
nor gate_2461(G1322,G1320,G1321);
nor gate_2462(G1325,G1323,G1324);
not gate_2463(G5392,G5388);
or gate_2464(G1790,G1708,G1789);
or gate_2465(G1982,G1941,G1981);
nand gate_2466(G1985,G5820,G5823);
nand gate_2467(G1988,G5828,G5831);
nand gate_2468(G1992,G5836,G5839);
nand gate_2469(G1995,G5844,G5847);
nand gate_2470(G2001,G1999,G2000);
not gate_2471(G2491,G2487);
and gate_2472(G2508,G2420,G2472,G2436,G2409,G2454);
and gate_2473(G2522,G4526,G2472,G2436,G2454,G2420);
and gate_2474(G2526,G4526,G2472,G2436,G2454);
and gate_2475(G2529,G4526,G2472,G2454);
and gate_2476(G2531,G4526,G2472);
not gate_2477(G5944,G5940);
not gate_2478(G5952,G5948);
not gate_2479(G5960,G5956);
not gate_2480(G5968,G5964);
nand gate_2481(G2555,G5972,G5975);
not gate_2482(G5976,G5972);
nand gate_2483(G2559,G5980,G5983);
not gate_2484(G5984,G5980);
not gate_2485(G2753,G2749);
and gate_2486(G2771,G2742,G2701,G2676,G2655,G2643);
and gate_2487(G2791,G2742,G2676,G2655,G2701);
and gate_2488(G2797,G2742,G2676,G2701);
and gate_2489(G2807,G2742,G2701);
not gate_2490(G6114,G6110);
not gate_2491(G6172,G6168);
not gate_2492(G6250,G6246);
not gate_2493(G6260,G6256);
not gate_2494(G6346,G6342);
not gate_2495(G6356,G6352);
not gate_2496(G3127,G3123);
and gate_2497(G3156,G3123,G3136);
or gate_2498(G3259,G3223,G3258);
and gate_2499(G3466,G3431,G3446);
not gate_2500(G6646,G6642);
not gate_2501(G6654,G6650);
not gate_2502(G6662,G6658);
not gate_2503(G6670,G6666);
nand gate_2504(G3483,G6674,G6677);
not gate_2505(G6678,G6674);
nand gate_2506(G3487,G6682,G6685);
not gate_2507(G6686,G6682);
not gate_2508(G3582,G3579);
not gate_2509(G3586,G3583);
not gate_2510(G3590,G3587);
not gate_2511(G3594,G3591);
nor gate_2512(G3597,G3595,G3596);
nor gate_2513(G3600,G3598,G3599);
and gate_2514(G3602,G3536,G3527,G3579);
and gate_2515(G3605,G3540,G3531,G3583);
and gate_2516(G3608,G3559,G3550,G3587);
and gate_2517(G3611,G3563,G3554,G3591);
not gate_2518(G4023,G4020);
not gate_2519(G6982,G6978);
not gate_2520(G7040,G7036);
not gate_2521(G7118,G7114);
not gate_2522(G7128,G7124);
and gate_2523(G4089,G4004,G4020);
not gate_2524(G4250,G4247);
not gate_2525(G4254,G4251);
not gate_2526(G4258,G4255);
not gate_2527(G4262,G4259);
and gate_2528(G4272,G4189,G4180,G4247);
and gate_2529(G4275,G4193,G4184,G4251);
and gate_2530(G4278,G4212,G4203,G4255);
and gate_2531(G4281,G4216,G4207,G4259);
nor gate_2532(G4285,G4283,G4284);
nor gate_2533(G4288,G4286,G4287);
not gate_2534(G4360,G4356);
nand gate_2535(G4380,G4369,G89);
and gate_2536(G4386,G4356,G4369);
not gate_2537(G7442,G7438);
not gate_2538(G4609,G4606);
not gate_2539(G4613,G4610);
not gate_2540(G4617,G4614);
not gate_2541(G4621,G4618);
nor gate_2542(G4624,G4622,G4623);
nor gate_2543(G4627,G4625,G4626);
and gate_2544(G4629,G4563,G4554,G4606);
and gate_2545(G4632,G4567,G4558,G4610);
and gate_2546(G4635,G4586,G4577,G4614);
and gate_2547(G4638,G4590,G4581,G4618);
buf gate_2548(G4836,G2472);
nand gate_2549(G4949,G4947,G4948);
nand gate_2550(G4990,G4988,G4989);
nand gate_2551(G5020,G5011,G5018);
nand gate_2552(G5108,G5099,G5106);
nand gate_2553(G5590,G5581,G5588);
nand gate_2554(G5678,G5669,G5676);
not gate_2555(G6084,G6080);
not gate_2556(G6094,G6090);
not gate_2557(G6104,G6100);
not gate_2558(G6142,G6138);
not gate_2559(G6152,G6148);
not gate_2560(G6162,G6158);
buf gate_2561(G6206,G2742);
not gate_2562(G6220,G6216);
not gate_2563(G6230,G6226);
not gate_2564(G6240,G6236);
not gate_2565(G6328,G6324);
buf gate_2566(G6294,G2742);
not gate_2567(G6308,G6304);
not gate_2568(G6318,G6314);
nand gate_2569(G6362,G6360,G6361);
nand gate_2570(G6840,G6817,G6818);
nand gate_2571(G6848,G6827,G6828);
not gate_2572(G6952,G6948);
not gate_2573(G6962,G6958);
not gate_2574(G6972,G6968);
not gate_2575(G7010,G7006);
not gate_2576(G7020,G7016);
not gate_2577(G7030,G7026);
not gate_2578(G7078,G7074);
not gate_2579(G7088,G7084);
not gate_2580(G7098,G7094);
not gate_2581(G7108,G7104);
not gate_2582(G7196,G7192);
not gate_2583(G7166,G7162);
not gate_2584(G7176,G7172);
not gate_2585(G7186,G7182);
nand gate_2586(G7448,G7446,G7447);
nand gate_2587(G7458,G7456,G7457);
and gate_2588(G254,G3046,G3249);
and gate_2589(G260,G3046,G3249);
nand gate_2590(G1987,G1985,G1986);
nand gate_2591(G1994,G1992,G1993);
not gate_2592(G2002,G2001);
and gate_2593(G962,G933,G924);
and gate_2594(G1751,G1730,G1721);
nand gate_2595(G1990,G1988,G1989);
nand gate_2596(G1997,G1995,G1996);
not gate_2597(G2499,G2495);
and gate_2598(G2536,G2515,G2487);
not gate_2599(G5943,G5937);
nand gate_2600(G2542,G5937,G5944);
not gate_2601(G5951,G5945);
nand gate_2602(G2545,G5945,G5952);
not gate_2603(G5959,G5953);
nand gate_2604(G2549,G5953,G5960);
not gate_2605(G5967,G5961);
nand gate_2606(G2552,G5961,G5968);
nand gate_2607(G2556,G5969,G5976);
nand gate_2608(G2560,G5977,G5984);
not gate_2609(G2761,G2757);
not gate_2610(G2784,G2780);
and gate_2611(G2853,G2749,G2780);
not gate_2612(G3135,G3131);
not gate_2613(G3146,G3143);
and gate_2614(G3163,G3123,G3143);
and gate_2615(G3467,G3453,G3431);
not gate_2616(G6645,G6639);
nand gate_2617(G3470,G6639,G6646);
not gate_2618(G6653,G6647);
nand gate_2619(G3473,G6647,G6654);
not gate_2620(G6661,G6655);
nand gate_2621(G3477,G6655,G6662);
not gate_2622(G6669,G6663);
nand gate_2623(G3480,G6663,G6670);
nand gate_2624(G3484,G6671,G6678);
nand gate_2625(G3488,G6679,G6686);
and gate_2626(G3601,G3531,G3536,G3582);
and gate_2627(G3604,G3527,G3540,G3586);
and gate_2628(G3607,G3554,G3559,G3590);
and gate_2629(G3610,G3550,G3563,G3594);
not gate_2630(G4032,G4028);
and gate_2631(G4090,G4004,G4028);
and gate_2632(G4271,G4184,G4189,G4250);
and gate_2633(G4274,G4180,G4193,G4254);
and gate_2634(G4277,G4207,G4212,G4258);
and gate_2635(G4280,G4203,G4216,G4262);
not gate_2636(G4368,G4364);
not gate_2637(G4379,G4376);
and gate_2638(G4387,G4356,G4376);
and gate_2639(G4628,G4558,G4563,G4609);
and gate_2640(G4631,G4554,G4567,G4613);
and gate_2641(G4634,G4581,G4586,G4617);
and gate_2642(G4637,G4577,G4590,G4621);
or gate_2643(G4841,G2431,G2518,G2519,G2520,G2522);
or gate_2644(G4849,G2448,G2523,G2524,G2526);
or gate_2645(G4857,G2465,G2527,G2529);
or gate_2646(G4865,G2481,G2531);
nand gate_2647(G5021,G5019,G5020);
not gate_2648(G5028,G5024);
nand gate_2649(G5109,G5107,G5108);
not gate_2650(G5116,G5112);
nand gate_2651(G5369,G1313,G1310);
nand gate_2652(G5377,G1319,G1316);
nand gate_2653(G5385,G1325,G1322);
not gate_2654(G5472,G5468);
nand gate_2655(G5473,G5468,G5471);
not gate_2656(G5530,G5526);
nand gate_2657(G5531,G5526,G5529);
nand gate_2658(G5591,G5589,G5590);
not gate_2659(G5598,G5594);
nand gate_2660(G5679,G5677,G5678);
not gate_2661(G5686,G5682);
or gate_2662(G6060,G2768,G2804);
not gate_2663(G6074,G6070);
not gate_2664(G6118,G2768);
not gate_2665(G6132,G6128);
or gate_2666(G6176,G2693,G2795,G2796,G2797);
or gate_2667(G6186,G2801,G2807);
or gate_2668(G6196,G2670,G2788,G2789,G2790,G2791);
not gate_2669(G6268,G6264);
nand gate_2670(G6269,G6264,G6267);
not gate_2671(G6274,G2801);
not gate_2672(G6288,G6284);
nand gate_2673(G6337,G4288,G4285);
nand gate_2674(G6829,G3600,G3597);
or gate_2675(G6928,G4017,G4051);
not gate_2676(G6942,G6938);
not gate_2677(G6986,G4017);
not gate_2678(G7000,G6996);
not gate_2679(G7048,G7044);
nand gate_2680(G7049,G7044,G7047);
or gate_2681(G7054,G4048,G4052);
not gate_2682(G7068,G7064);
not gate_2683(G7136,G7132);
nand gate_2684(G7137,G7132,G7135);
not gate_2685(G7142,G4048);
not gate_2686(G7156,G7152);
nand gate_2687(G7433,G4627,G4624);
and gate_2688(G242,G1982,G1146);
nand gate_2689(G3151,G3135,G3127);
and gate_2690(G257,G89,G4386,G3156,G3035,G3249);
and gate_2691(G263,G89,G4386,G3156,G3035,G3249);
and gate_2692(G266,G1790,G997);
not gate_2693(G1991,G1990);
not gate_2694(G1998,G1997);
nand gate_2695(G3489,G3487,G3488);
nand gate_2696(G371,G4836,G4839);
not gate_2697(G4840,G4836);
nand gate_2698(G2561,G2559,G2560);
and gate_2699(G2532,G2487,G2508);
or gate_2700(G2537,G2495,G2536);
nand gate_2701(G2541,G5940,G5943);
nand gate_2702(G2544,G5948,G5951);
nand gate_2703(G2548,G5956,G5959);
nand gate_2704(G2551,G5964,G5967);
nand gate_2705(G2557,G2555,G2556);
and gate_2706(G2563,G2508,G4526);
nand gate_2707(G2577,G2499,G2491);
not gate_2708(G2775,G2771);
nand gate_2709(G2806,G2771,G4526);
nand gate_2710(G2808,G2761,G2753);
and gate_2711(G2852,G2749,G2771);
or gate_2712(G2854,G2757,G2853);
not gate_2713(G6366,G6362);
nand gate_2714(G4381,G4368,G4360);
or gate_2715(G3164,G3131,G3163);
and gate_2716(G3241,G89,G4386,G3156,G3035);
or gate_2717(G3468,G3437,G3467);
nand gate_2718(G3469,G6642,G6645);
nand gate_2719(G3472,G6650,G6653);
nand gate_2720(G3476,G6658,G6661);
nand gate_2721(G3479,G6666,G6669);
nand gate_2722(G3485,G3483,G3484);
nor gate_2723(G3603,G3601,G3602);
nor gate_2724(G3606,G3604,G3605);
nor gate_2725(G3609,G3607,G3608);
nor gate_2726(G3612,G3610,G3611);
not gate_2727(G6844,G6840);
not gate_2728(G6852,G6848);
or gate_2729(G4091,G4010,G4090);
nor gate_2730(G4273,G4271,G4272);
nor gate_2731(G4276,G4274,G4275);
nor gate_2732(G4279,G4277,G4278);
nor gate_2733(G4282,G4280,G4281);
and gate_2734(G4382,G4379,G4380);
or gate_2735(G4388,G4364,G4387);
not gate_2736(G7452,G7448);
not gate_2737(G7462,G7458);
nor gate_2738(G4630,G4628,G4629);
nor gate_2739(G4633,G4631,G4632);
nor gate_2740(G4636,G4634,G4635);
nor gate_2741(G4639,G4637,G4638);
not gate_2742(G4955,G4949);
nand gate_2743(G4958,G4949,G4956);
not gate_2744(G4996,G4990);
nand gate_2745(G4999,G4990,G4997);
nand gate_2746(G5474,G5465,G5472);
nand gate_2747(G5532,G5523,G5530);
not gate_2748(G6210,G6206);
nand gate_2749(G6270,G6261,G6268);
not gate_2750(G6298,G6294);
nand gate_2751(G7050,G7041,G7048);
nand gate_2752(G7138,G7129,G7136);
nand gate_2753(G3471,G3469,G3470);
nand gate_2754(G3478,G3476,G3477);
not gate_2755(G3486,G3485);
nand gate_2756(G372,G4833,G4840);
nand gate_2757(G2543,G2541,G2542);
nand gate_2758(G2550,G2548,G2549);
not gate_2759(G2558,G2557);
not gate_2760(G4847,G4841);
nand gate_2761(G387,G4841,G4848);
not gate_2762(G4855,G4849);
nand gate_2763(G390,G4849,G4856);
not gate_2764(G4863,G4857);
nand gate_2765(G393,G4857,G4864);
not gate_2766(G4871,G4865);
nand gate_2767(G396,G4865,G4872);
not gate_2768(G965,G962);
not gate_2769(G5375,G5369);
nand gate_2770(G1327,G5369,G5376);
not gate_2771(G5383,G5377);
nand gate_2772(G1330,G5377,G5384);
not gate_2773(G5391,G5385);
nand gate_2774(G1333,G5385,G5392);
not gate_2775(G1754,G1751);
nand gate_2776(G2546,G2544,G2545);
nand gate_2777(G2553,G2551,G2552);
or gate_2778(G2564,G2515,G2563);
and gate_2779(G2809,G2784,G2806);
and gate_2780(G2813,G2784,G2775);
not gate_2781(G6345,G6337);
nand gate_2782(G2860,G6337,G6346);
nand gate_2783(G3474,G3472,G3473);
nand gate_2784(G3481,G3479,G3480);
not gate_2785(G6835,G6829);
nand gate_2786(G3614,G6829,G6836);
and gate_2787(G4053,G4032,G4023);
not gate_2788(G7441,G7433);
nand gate_2789(G4516,G7433,G7442);
nand gate_2790(G4957,G4952,G4955);
nand gate_2791(G4998,G4993,G4996);
not gate_2792(G5027,G5021);
nand gate_2793(G5030,G5021,G5028);
not gate_2794(G5115,G5109);
nand gate_2795(G5118,G5109,G5116);
nand gate_2796(G5475,G5473,G5474);
nand gate_2797(G5533,G5531,G5532);
not gate_2798(G5597,G5591);
nand gate_2799(G5600,G5591,G5598);
not gate_2800(G5685,G5679);
nand gate_2801(G5688,G5679,G5686);
not gate_2802(G6064,G6060);
nand gate_2803(G6065,G6060,G6063);
not gate_2804(G6122,G6118);
nand gate_2805(G6123,G6118,G6121);
not gate_2806(G6180,G6176);
nand gate_2807(G6181,G6176,G6179);
not gate_2808(G6190,G6186);
not gate_2809(G6200,G6196);
nand gate_2810(G6271,G6269,G6270);
not gate_2811(G6278,G6274);
nand gate_2812(G6347,G4276,G4273);
nand gate_2813(G6357,G4282,G4279);
nand gate_2814(G6837,G3606,G3603);
nand gate_2815(G6845,G3612,G3609);
not gate_2816(G6932,G6928);
nand gate_2817(G6933,G6928,G6931);
not gate_2818(G6990,G6986);
nand gate_2819(G6991,G6986,G6989);
nand gate_2820(G7051,G7049,G7050);
not gate_2821(G7058,G7054);
nand gate_2822(G7139,G7137,G7138);
not gate_2823(G7146,G7142);
nand gate_2824(G7443,G4639,G4636);
nand gate_2825(G7453,G4633,G4630);
and gate_2826(G243,G3468,G1974,G1146);
and gate_2827(G244,G2537,G3466,G1974,G1146);
and gate_2828(G245,G4526,G2532,G3466,G1974,G1146);
and gate_2829(G255,G3164,G3035,G3249);
and gate_2830(G256,G4388,G3156,G3035,G3249);
and gate_2831(G261,G3164,G3035,G3249);
and gate_2832(G262,G4388,G3156,G3035,G3249);
and gate_2833(G267,G4091,G1788,G997);
and gate_2834(G268,G2854,G4089,G1788,G997);
and gate_2835(G269,G4526,G2852,G4089,G1788,G997);
not gate_2836(G3475,G3474);
not gate_2837(G3482,G3481);
nand gate_2838(G373,G371,G372);
not gate_2839(G2547,G2546);
not gate_2840(G2554,G2553);
nand gate_2841(G386,G4844,G4847);
nand gate_2842(G389,G4852,G4855);
nand gate_2843(G392,G4860,G4863);
nand gate_2844(G395,G4868,G4871);
nand gate_2845(G1326,G5372,G5375);
nand gate_2846(G1329,G5380,G5383);
nand gate_2847(G1332,G5388,G5391);
and gate_2848(G1436,G4091,G1788);
and gate_2849(G1440,G2854,G4089,G1788);
and gate_2850(G1445,G4526,G2852,G4089,G1788);
and gate_2851(G1450,G2854,G4089);
and gate_2852(G1454,G4526,G2852,G4089);
nand gate_2853(G2859,G6342,G6345);
not gate_2854(G4385,G4382);
and gate_2855(G3148,G4382,G4364);
and gate_2856(G3239,G3164,G3035);
and gate_2857(G3240,G4388,G3156,G3035);
and gate_2858(G3265,G3468,G1974);
and gate_2859(G3267,G2537,G3466,G1974);
and gate_2860(G3270,G4526,G2532,G3466,G1974);
and gate_2861(G3274,G2537,G3466);
and gate_2862(G3277,G4526,G2532,G3466);
nand gate_2863(G3613,G6832,G6835);
nand gate_2864(G4515,G7438,G7441);
nand gate_2865(G4959,G4957,G4958);
nand gate_2866(G5000,G4998,G4999);
nand gate_2867(G5029,G5024,G5027);
nand gate_2868(G5117,G5112,G5115);
nand gate_2869(G5599,G5594,G5597);
nand gate_2870(G5687,G5682,G5685);
nand gate_2871(G6066,G6057,G6064);
nand gate_2872(G6124,G6115,G6122);
nand gate_2873(G6182,G6173,G6180);
nand gate_2874(G6934,G6925,G6932);
nand gate_2875(G6992,G6983,G6990);
or gate_2876(G246,G241,G242,G243,G244,G245);
or gate_2877(G258,G3259,G254,G255,G256,G257);
or gate_2878(G264,G3259,G260,G261,G262,G263);
or gate_2879(G270,G265,G266,G267,G268,G269);
and gate_2880(G375,G2564,G2543);
and gate_2881(G378,G2564,G2550);
and gate_2882(G381,G2564,G2558);
and gate_2883(G384,G2564,G2406);
nand gate_2884(G388,G386,G387);
nand gate_2885(G391,G389,G390);
nand gate_2886(G394,G392,G393);
nand gate_2887(G397,G395,G396);
nand gate_2888(G1328,G1326,G1327);
nand gate_2889(G1331,G1329,G1330);
nand gate_2890(G1334,G1332,G1333);
or gate_2891(G1447,G1790,G1436,G1440,G1445);
or gate_2892(G1766,G4091,G1450,G1454);
not gate_2893(G2571,G2564);
and gate_2894(G2579,G2577,G2564);
not gate_2895(G2812,G2809);
not gate_2896(G2816,G2813);
and gate_2897(G2851,G2809,G2757);
nand gate_2898(G2861,G2859,G2860);
not gate_2899(G6355,G6347);
nand gate_2900(G2863,G6347,G6356);
not gate_2901(G6365,G6357);
nand gate_2902(G2866,G6357,G6366);
and gate_2903(G3147,G4381,G4385);
or gate_2904(G3242,G3046,G3239,G3240,G3241);
or gate_2905(G3271,G1982,G3265,G3267,G3270);
or gate_2906(G3279,G3468,G3274,G3277);
nand gate_2907(G3615,G3613,G3614);
not gate_2908(G6843,G6837);
nand gate_2909(G3617,G6837,G6844);
not gate_2910(G6851,G6845);
nand gate_2911(G3620,G6845,G6852);
not gate_2912(G4056,G4053);
nand gate_2913(G4517,G4515,G4516);
not gate_2914(G7451,G7443);
nand gate_2915(G4519,G7443,G7452);
not gate_2916(G7461,G7453);
nand gate_2917(G4522,G7453,G7462);
nand gate_2918(G5031,G5029,G5030);
nand gate_2919(G5119,G5117,G5118);
not gate_2920(G5481,G5475);
nand gate_2921(G5484,G5475,G5482);
not gate_2922(G5539,G5533);
nand gate_2923(G5542,G5533,G5540);
nand gate_2924(G5601,G5599,G5600);
nand gate_2925(G5689,G5687,G5688);
nand gate_2926(G6067,G6065,G6066);
nand gate_2927(G6125,G6123,G6124);
nand gate_2928(G6183,G6181,G6182);
not gate_2929(G6277,G6271);
nand gate_2930(G6280,G6271,G6278);
nand gate_2931(G6935,G6933,G6934);
nand gate_2932(G6993,G6991,G6992);
not gate_2933(G7057,G7051);
nand gate_2934(G7060,G7051,G7058);
not gate_2935(G7145,G7139);
nand gate_2936(G7148,G7139,G7146);
nand gate_2937(G4968,G4959,G4966);
nand gate_2938(G5009,G5000,G5007);
and gate_2939(G2850,G2808,G2812);
nand gate_2940(G2862,G6352,G6355);
nand gate_2941(G2865,G6362,G6365);
or gate_2942(G3149,G3147,G3148);
nand gate_2943(G3243,G3228,G3242);
nand gate_2944(G3616,G6840,G6843);
nand gate_2945(G3619,G6848,G6851);
nand gate_2946(G4518,G7448,G7451);
nand gate_2947(G4521,G7458,G7461);
not gate_2948(G4965,G4959);
not gate_2949(G5006,G5000);
nand gate_2950(G5483,G5478,G5481);
nand gate_2951(G5541,G5536,G5539);
nand gate_2952(G6279,G6274,G6277);
nand gate_2953(G7059,G7054,G7057);
nand gate_2954(G7147,G7142,G7145);
and gate_2955(G374,G2547,G2571);
and gate_2956(G377,G2554,G2571);
and gate_2957(G380,G2561,G2571);
and gate_2958(G383,G2400,G2571);
nand gate_2959(G955,G920,G1447);
nand gate_2960(G4967,G4962,G4965);
nand gate_2961(G5008,G5003,G5006);
buf gate_2962(G975,G1447);
and gate_2963(G1136,G3271,G1093,G1055,G1074,G1038);
and gate_2964(G1140,G3271,G1093,G1055,G1074);
and gate_2965(G1143,G3271,G1093,G1074);
and gate_2966(G1145,G3271,G1093);
and gate_2967(G1160,G1122,G3271);
not gate_2968(G1771,G1766);
and gate_2969(G1964,G3279,G1921,G1885,G1903,G1869);
and gate_2970(G1968,G3279,G1921,G1885,G1903);
and gate_2971(G1971,G3279,G1921,G1903);
and gate_2972(G1973,G3279,G1921);
and gate_2973(G2007,G1950,G3279);
and gate_2974(G2578,G2495,G2571);
nand gate_2975(G2864,G2862,G2863);
nand gate_2976(G2867,G2865,G2866);
nand gate_2977(G3150,G3136,G3149);
and gate_2978(G3245,G3238,G3243);
nand gate_2979(G3618,G3616,G3617);
nand gate_2980(G3621,G3619,G3620);
or gate_2981(G4067,G2850,G2851);
nand gate_2982(G4520,G4518,G4519);
nand gate_2983(G4523,G4521,G4522);
buf gate_2984(G4713,G3279);
buf gate_2985(G4753,G3271);
not gate_2986(G5037,G5031);
nand gate_2987(G5040,G5031,G5038);
not gate_2988(G5125,G5119);
nand gate_2989(G5128,G5119,G5126);
nand gate_2990(G5485,G5483,G5484);
nand gate_2991(G5543,G5541,G5542);
not gate_2992(G5607,G5601);
nand gate_2993(G5610,G5601,G5608);
not gate_2994(G5695,G5689);
nand gate_2995(G5698,G5689,G5696);
not gate_2996(G6073,G6067);
nand gate_2997(G6076,G6067,G6074);
not gate_2998(G6131,G6125);
nand gate_2999(G6134,G6125,G6132);
not gate_3000(G6189,G6183);
nand gate_3001(G6192,G6183,G6190);
nand gate_3002(G6281,G6279,G6280);
not gate_3003(G6941,G6935);
nand gate_3004(G6944,G6935,G6942);
not gate_3005(G6999,G6993);
nand gate_3006(G7002,G6993,G7000);
nand gate_3007(G7061,G7059,G7060);
nand gate_3008(G7149,G7147,G7148);
or gate_3009(G376,G374,G375);
or gate_3010(G379,G377,G378);
or gate_3011(G382,G380,G381);
or gate_3012(G385,G383,G384);
and gate_3013(G958,G933,G955);
nand gate_3014(G967,G4967,G4968);
nand gate_3015(G971,G5008,G5009);
or gate_3016(G1161,G1129,G1160);
or gate_3017(G2008,G1957,G2007);
or gate_3018(G2580,G2578,G2579);
and gate_3019(G2868,G1331,G2861,G2864,G2867);
and gate_3020(G3152,G3146,G3150);
and gate_3021(G4443,G1328,G1334,G3618,G3621);
and gate_3022(G4524,G3615,G4517,G4520,G4523);
or gate_3023(G4721,G1880,G1960,G1961,G1962,G1964);
or gate_3024(G4729,G1897,G1965,G1966,G1968);
or gate_3025(G4737,G1914,G1969,G1971);
or gate_3026(G4745,G1929,G1973);
or gate_3027(G4761,G1050,G1132,G1133,G1134,G1136);
or gate_3028(G4769,G1068,G1137,G1138,G1140);
or gate_3029(G4777,G1086,G1141,G1143);
or gate_3030(G4785,G1102,G1145);
nand gate_3031(G5039,G5034,G5037);
nand gate_3032(G5127,G5122,G5125);
nand gate_3033(G5609,G5604,G5607);
nand gate_3034(G5697,G5692,G5695);
nand gate_3035(G6075,G6070,G6073);
nand gate_3036(G6133,G6128,G6131);
nand gate_3037(G6191,G6186,G6189);
nand gate_3038(G6943,G6938,G6941);
nand gate_3039(G7001,G6996,G6999);
not gate_3040(G3248,G3245);
and gate_3041(G248,G3245,G3223);
not gate_3042(G4719,G4713);
nand gate_3043(G294,G4713,G4720);
not gate_3044(G4759,G4753);
nand gate_3045(G323,G4753,G4760);
not gate_3046(G980,G975);
not gate_3047(G4072,G4067);
nand gate_3048(G5041,G5039,G5040);
nand gate_3049(G5129,G5127,G5128);
not gate_3050(G5491,G5485);
nand gate_3051(G5494,G5485,G5492);
not gate_3052(G5549,G5543);
nand gate_3053(G5552,G5543,G5550);
nand gate_3054(G5611,G5609,G5610);
nand gate_3055(G5699,G5697,G5698);
nand gate_3056(G6077,G6075,G6076);
nand gate_3057(G6135,G6133,G6134);
nand gate_3058(G6193,G6191,G6192);
not gate_3059(G6287,G6281);
nand gate_3060(G6290,G6281,G6288);
nand gate_3061(G6945,G6943,G6944);
nand gate_3062(G7003,G7001,G7002);
not gate_3063(G7067,G7061);
nand gate_3064(G7070,G7061,G7068);
not gate_3065(G7155,G7149);
nand gate_3066(G7158,G7149,G7156);
and gate_3067(G247,G3244,G3248);
not gate_3068(G3155,G3152);
and gate_3069(G251,G3152,G3131);
and gate_3070(G272,G1176,G1161);
not gate_3071(G961,G958);
and gate_3072(G275,G958,G908);
nand gate_3073(G293,G4716,G4719);
and gate_3074(G297,G2008,G1987);
and gate_3075(G300,G2008,G1994);
and gate_3076(G303,G2008,G2002);
and gate_3077(G306,G2008,G1856);
not gate_3078(G4727,G4721);
nand gate_3079(G309,G4721,G4728);
not gate_3080(G4735,G4729);
nand gate_3081(G312,G4729,G4736);
not gate_3082(G4743,G4737);
nand gate_3083(G315,G4737,G4744);
not gate_3084(G4751,G4745);
nand gate_3085(G318,G4745,G4752);
nand gate_3086(G322,G4756,G4759);
not gate_3087(G4767,G4761);
nand gate_3088(G326,G4761,G4768);
not gate_3089(G4775,G4769);
nand gate_3090(G329,G4769,G4776);
not gate_3091(G4783,G4777);
nand gate_3092(G332,G4777,G4784);
not gate_3093(G4791,G4785);
nand gate_3094(G335,G4785,G4792);
not gate_3095(G412,G4443);
not gate_3096(G414,G4524);
not gate_3097(G416,G2868);
and gate_3098(G2881,G4443,G4524,G2868);
and gate_3099(G993,G971,G962,G975);
and gate_3100(G994,G967,G965,G975);
not gate_3101(G1166,G1161);
and gate_3102(G1171,G1161,G1155);
and gate_3103(G1174,G1161,G1023);
not gate_3104(G2014,G2008);
and gate_3105(G3459,G2580,G3417,G3381,G3399,G3365);
and gate_3106(G3462,G2580,G3417,G3381,G3399);
and gate_3107(G3464,G2580,G3417,G3399);
and gate_3108(G3465,G2580,G3417);
and gate_3109(G3490,G3446,G2580);
buf gate_3110(G4793,G2580);
nand gate_3111(G5493,G5488,G5491);
nand gate_3112(G5551,G5546,G5549);
nand gate_3113(G6289,G6284,G6287);
nand gate_3114(G7069,G7064,G7067);
nand gate_3115(G7157,G7152,G7155);
or gate_3116(G249,G247,G248);
and gate_3117(G250,G3151,G3155);
and gate_3118(G274,G957,G961);
nand gate_3119(G295,G293,G294);
nand gate_3120(G308,G4724,G4727);
nand gate_3121(G311,G4732,G4735);
nand gate_3122(G314,G4740,G4743);
nand gate_3123(G317,G4748,G4751);
nand gate_3124(G324,G322,G323);
nand gate_3125(G325,G4764,G4767);
nand gate_3126(G328,G4772,G4775);
nand gate_3127(G331,G4780,G4783);
nand gate_3128(G334,G4788,G4791);
and gate_3129(G417,G2876,G2878,G2881);
and gate_3130(G991,G971,G933,G980);
and gate_3131(G992,G967,G929,G980);
or gate_3132(G3491,G3453,G3490);
or gate_3133(G4801,G3376,G3456,G3457,G3458,G3459);
or gate_3134(G4809,G3393,G3460,G3461,G3462);
or gate_3135(G4817,G3410,G3463,G3464);
or gate_3136(G4825,G3425,G3465);
not gate_3137(G5047,G5041);
nand gate_3138(G5050,G5041,G5048);
not gate_3139(G5135,G5129);
nand gate_3140(G5138,G5129,G5136);
nand gate_3141(G5495,G5493,G5494);
nand gate_3142(G5553,G5551,G5552);
not gate_3143(G5617,G5611);
nand gate_3144(G5620,G5611,G5618);
not gate_3145(G5705,G5699);
nand gate_3146(G5708,G5699,G5706);
not gate_3147(G6083,G6077);
nand gate_3148(G6086,G6077,G6084);
not gate_3149(G6141,G6135);
nand gate_3150(G6144,G6135,G6142);
not gate_3151(G6199,G6193);
nand gate_3152(G6202,G6193,G6200);
nand gate_3153(G6291,G6289,G6290);
not gate_3154(G6951,G6945);
nand gate_3155(G6954,G6945,G6952);
not gate_3156(G7009,G7003);
nand gate_3157(G7012,G7003,G7010);
nand gate_3158(G7071,G7069,G7070);
nand gate_3159(G7159,G7157,G7158);
or gate_3160(G252,G250,G251);
and gate_3161(G271,G1117,G1166);
or gate_3162(G276,G274,G275);
and gate_3163(G296,G1991,G2014);
and gate_3164(G299,G1998,G2014);
and gate_3165(G302,G2005,G2014);
and gate_3166(G305,G1850,G2014);
nand gate_3167(G310,G308,G309);
nand gate_3168(G313,G311,G312);
nand gate_3169(G316,G314,G315);
nand gate_3170(G319,G317,G318);
nand gate_3171(G327,G325,G326);
nand gate_3172(G330,G328,G329);
nand gate_3173(G333,G331,G332);
nand gate_3174(G336,G334,G335);
not gate_3175(G4799,G4793);
nand gate_3176(G343,G4793,G4800);
not gate_3177(G418,G417);
and gate_3178(G1170,G1158,G1166);
and gate_3179(G1173,G1019,G1166);
nand gate_3180(G5049,G5044,G5047);
nand gate_3181(G5137,G5132,G5135);
or gate_3182(G5167,G991,G992,G993,G994);
nand gate_3183(G5619,G5614,G5617);
nand gate_3184(G5707,G5702,G5705);
nand gate_3185(G6085,G6080,G6083);
nand gate_3186(G6143,G6138,G6141);
nand gate_3187(G6201,G6196,G6199);
nand gate_3188(G6953,G6948,G6951);
nand gate_3189(G7011,G7006,G7009);
or gate_3190(G273,G271,G272);
or gate_3191(G298,G296,G297);
or gate_3192(G301,G299,G300);
or gate_3193(G304,G302,G303);
or gate_3194(G307,G305,G306);
nand gate_3195(G342,G4796,G4799);
and gate_3196(G346,G3491,G3471);
and gate_3197(G349,G3491,G3478);
and gate_3198(G352,G3491,G3486);
and gate_3199(G355,G3491,G3350);
not gate_3200(G4807,G4801);
nand gate_3201(G358,G4801,G4808);
not gate_3202(G4815,G4809);
nand gate_3203(G361,G4809,G4816);
not gate_3204(G4823,G4817);
nand gate_3205(G364,G4817,G4824);
not gate_3206(G4831,G4825);
nand gate_3207(G367,G4825,G4832);
or gate_3208(G1172,G1170,G1171);
or gate_3209(G1175,G1173,G1174);
not gate_3210(G3497,G3491);
nand gate_3211(G5051,G5049,G5050);
nand gate_3212(G5139,G5137,G5138);
not gate_3213(G5501,G5495);
nand gate_3214(G5504,G5495,G5502);
not gate_3215(G5559,G5553);
nand gate_3216(G5562,G5553,G5560);
nand gate_3217(G5621,G5619,G5620);
nand gate_3218(G5709,G5707,G5708);
nand gate_3219(G6087,G6085,G6086);
nand gate_3220(G6145,G6143,G6144);
nand gate_3221(G6203,G6201,G6202);
not gate_3222(G6297,G6291);
nand gate_3223(G6300,G6291,G6298);
nand gate_3224(G6955,G6953,G6954);
nand gate_3225(G7013,G7011,G7012);
not gate_3226(G7077,G7071);
nand gate_3227(G7080,G7071,G7078);
not gate_3228(G7165,G7159);
nand gate_3229(G7168,G7159,G7166);
nand gate_3230(G344,G342,G343);
nand gate_3231(G357,G4804,G4807);
nand gate_3232(G360,G4812,G4815);
nand gate_3233(G363,G4820,G4823);
nand gate_3234(G366,G4828,G4831);
not gate_3235(G5173,G5167);
buf gate_3236(G422,G1172);
buf gate_3237(G469,G1172);
buf gate_3238(G419,G1175);
buf gate_3239(G471,G1175);
nand gate_3240(G5503,G5498,G5501);
nand gate_3241(G5561,G5556,G5559);
nand gate_3242(G6299,G6294,G6297);
nand gate_3243(G7079,G7074,G7077);
nand gate_3244(G7167,G7162,G7165);
and gate_3245(G345,G3475,G3497);
and gate_3246(G348,G3482,G3497);
and gate_3247(G351,G3489,G3497);
and gate_3248(G354,G3344,G3497);
nand gate_3249(G359,G357,G358);
nand gate_3250(G362,G360,G361);
nand gate_3251(G365,G363,G364);
nand gate_3252(G368,G366,G367);
not gate_3253(G5057,G5051);
nand gate_3254(G5060,G5051,G5058);
not gate_3255(G5145,G5139);
nand gate_3256(G5148,G5139,G5146);
nand gate_3257(G5505,G5503,G5504);
nand gate_3258(G5563,G5561,G5562);
not gate_3259(G5627,G5621);
nand gate_3260(G5630,G5621,G5628);
not gate_3261(G5715,G5709);
nand gate_3262(G5718,G5709,G5716);
not gate_3263(G6093,G6087);
nand gate_3264(G6096,G6087,G6094);
not gate_3265(G6151,G6145);
nand gate_3266(G6154,G6145,G6152);
not gate_3267(G6209,G6203);
nand gate_3268(G6212,G6203,G6210);
nand gate_3269(G6301,G6299,G6300);
not gate_3270(G6961,G6955);
nand gate_3271(G6964,G6955,G6962);
not gate_3272(G7019,G7013);
nand gate_3273(G7022,G7013,G7020);
nand gate_3274(G7081,G7079,G7080);
nand gate_3275(G7169,G7167,G7168);
or gate_3276(G347,G345,G346);
or gate_3277(G350,G348,G349);
or gate_3278(G353,G351,G352);
or gate_3279(G356,G354,G355);
nand gate_3280(G5059,G5054,G5057);
nand gate_3281(G5147,G5142,G5145);
nand gate_3282(G5629,G5624,G5627);
nand gate_3283(G5717,G5712,G5715);
nand gate_3284(G6095,G6090,G6093);
nand gate_3285(G6153,G6148,G6151);
nand gate_3286(G6211,G6206,G6209);
nand gate_3287(G6963,G6958,G6961);
nand gate_3288(G7021,G7016,G7019);
nand gate_3289(G5061,G5059,G5060);
nand gate_3290(G5149,G5147,G5148);
not gate_3291(G5511,G5505);
nand gate_3292(G5514,G5505,G5512);
not gate_3293(G5569,G5563);
nand gate_3294(G5572,G5563,G5570);
nand gate_3295(G5631,G5629,G5630);
nand gate_3296(G5719,G5717,G5718);
nand gate_3297(G6097,G6095,G6096);
nand gate_3298(G6155,G6153,G6154);
nand gate_3299(G6213,G6211,G6212);
not gate_3300(G6307,G6301);
nand gate_3301(G6310,G6301,G6308);
nand gate_3302(G6965,G6963,G6964);
nand gate_3303(G7023,G7021,G7022);
not gate_3304(G7087,G7081);
nand gate_3305(G7090,G7081,G7088);
not gate_3306(G7175,G7169);
nand gate_3307(G7178,G7169,G7176);
nand gate_3308(G5513,G5508,G5511);
nand gate_3309(G5571,G5566,G5569);
nand gate_3310(G6309,G6304,G6307);
nand gate_3311(G7089,G7084,G7087);
nand gate_3312(G7177,G7172,G7175);
not gate_3313(G5067,G5061);
nand gate_3314(G5070,G5061,G5068);
not gate_3315(G5155,G5149);
nand gate_3316(G5158,G5149,G5156);
nand gate_3317(G5515,G5513,G5514);
nand gate_3318(G5573,G5571,G5572);
not gate_3319(G5637,G5631);
nand gate_3320(G5640,G5631,G5638);
not gate_3321(G5725,G5719);
nand gate_3322(G5728,G5719,G5726);
not gate_3323(G6103,G6097);
nand gate_3324(G6106,G6097,G6104);
not gate_3325(G6161,G6155);
nand gate_3326(G6164,G6155,G6162);
not gate_3327(G6219,G6213);
nand gate_3328(G6222,G6213,G6220);
nand gate_3329(G6311,G6309,G6310);
not gate_3330(G6971,G6965);
nand gate_3331(G6974,G6965,G6972);
not gate_3332(G7029,G7023);
nand gate_3333(G7032,G7023,G7030);
nand gate_3334(G7091,G7089,G7090);
nand gate_3335(G7179,G7177,G7178);
nand gate_3336(G5069,G5064,G5067);
nand gate_3337(G5157,G5152,G5155);
nand gate_3338(G5639,G5634,G5637);
nand gate_3339(G5727,G5722,G5725);
nand gate_3340(G6105,G6100,G6103);
nand gate_3341(G6163,G6158,G6161);
nand gate_3342(G6221,G6216,G6219);
nand gate_3343(G6973,G6968,G6971);
nand gate_3344(G7031,G7026,G7029);
not gate_3345(G5521,G5515);
nand gate_3346(G1756,G5515,G5522);
not gate_3347(G5579,G5573);
nand gate_3348(G1761,G5573,G5580);
nand gate_3349(G5071,G5069,G5070);
nand gate_3350(G5159,G5157,G5158);
nand gate_3351(G5641,G5639,G5640);
nand gate_3352(G5729,G5727,G5728);
nand gate_3353(G6107,G6105,G6106);
nand gate_3354(G6165,G6163,G6164);
nand gate_3355(G6223,G6221,G6222);
not gate_3356(G6317,G6311);
nand gate_3357(G6320,G6311,G6318);
nand gate_3358(G6975,G6973,G6974);
nand gate_3359(G7033,G7031,G7032);
not gate_3360(G7097,G7091);
nand gate_3361(G7100,G7091,G7098);
not gate_3362(G7185,G7179);
nand gate_3363(G7188,G7179,G7186);
nand gate_3364(G1755,G5518,G5521);
nand gate_3365(G1760,G5576,G5579);
nand gate_3366(G6319,G6314,G6317);
nand gate_3367(G7099,G7094,G7097);
nand gate_3368(G7187,G7182,G7185);
nand gate_3369(G1757,G1755,G1756);
nand gate_3370(G1762,G1760,G1761);
not gate_3371(G6113,G6107);
nand gate_3372(G2818,G6107,G6114);
not gate_3373(G6171,G6165);
nand gate_3374(G2823,G6165,G6172);
not gate_3375(G6981,G6975);
nand gate_3376(G4058,G6975,G6982);
not gate_3377(G7039,G7033);
nand gate_3378(G4063,G7033,G7040);
not gate_3379(G5077,G5071);
nand gate_3380(G5080,G5071,G5078);
not gate_3381(G5165,G5159);
nand gate_3382(G5090,G5159,G5166);
not gate_3383(G5647,G5641);
nand gate_3384(G5650,G5641,G5648);
not gate_3385(G5735,G5729);
nand gate_3386(G5660,G5729,G5736);
not gate_3387(G6229,G6223);
nand gate_3388(G6232,G6223,G6230);
nand gate_3389(G6321,G6319,G6320);
nand gate_3390(G7101,G7099,G7100);
nand gate_3391(G7189,G7187,G7188);
nand gate_3392(G2817,G6110,G6113);
nand gate_3393(G2822,G6168,G6171);
nand gate_3394(G4057,G6978,G6981);
nand gate_3395(G4062,G7036,G7039);
nand gate_3396(G5079,G5074,G5077);
nand gate_3397(G5089,G5162,G5165);
nand gate_3398(G5649,G5644,G5647);
nand gate_3399(G5659,G5732,G5735);
nand gate_3400(G6231,G6226,G6229);
and gate_3401(G1782,G1762,G1730,G1771);
and gate_3402(G1783,G1757,G1726,G1771);
and gate_3403(G1784,G1762,G1751,G1766);
and gate_3404(G1785,G1757,G1754,G1766);
nand gate_3405(G2819,G2817,G2818);
nand gate_3406(G2824,G2822,G2823);
nand gate_3407(G4059,G4057,G4058);
nand gate_3408(G4064,G4062,G4063);
nand gate_3409(G5081,G5079,G5080);
nand gate_3410(G5091,G5089,G5090);
nand gate_3411(G5651,G5649,G5650);
nand gate_3412(G5661,G5659,G5660);
nand gate_3413(G6233,G6231,G6232);
not gate_3414(G6327,G6321);
nand gate_3415(G6252,G6321,G6328);
not gate_3416(G7107,G7101);
nand gate_3417(G7110,G7101,G7108);
not gate_3418(G7195,G7189);
nand gate_3419(G7120,G7189,G7196);
or gate_3420(G5737,G1782,G1783,G1784,G1785);
nand gate_3421(G6251,G6324,G6327);
nand gate_3422(G7109,G7104,G7107);
nand gate_3423(G7119,G7192,G7195);
not gate_3424(G5087,G5081);
nand gate_3425(G985,G5081,G5088);
not gate_3426(G5097,G5091);
nand gate_3427(G988,G5091,G5098);
not gate_3428(G5657,G5651);
nand gate_3429(G1776,G5651,G5658);
not gate_3430(G5667,G5661);
nand gate_3431(G1779,G5661,G5668);
and gate_3432(G2844,G2824,G2784,G2833);
and gate_3433(G2845,G2819,G2780,G2833);
and gate_3434(G2846,G2824,G2813,G2828);
and gate_3435(G2847,G2819,G2816,G2828);
and gate_3436(G4083,G4064,G4032,G4072);
and gate_3437(G4084,G4059,G4028,G4072);
and gate_3438(G4085,G4064,G4053,G4067);
and gate_3439(G4086,G4059,G4056,G4067);
not gate_3440(G6239,G6233);
nand gate_3441(G6242,G6233,G6240);
nand gate_3442(G6253,G6251,G6252);
nand gate_3443(G7111,G7109,G7110);
nand gate_3444(G7121,G7119,G7120);
nand gate_3445(G984,G5084,G5087);
nand gate_3446(G987,G5094,G5097);
nand gate_3447(G1775,G5654,G5657);
nand gate_3448(G1778,G5664,G5667);
not gate_3449(G5743,G5737);
nand gate_3450(G6241,G6236,G6239);
or gate_3451(G6329,G2844,G2845,G2846,G2847);
or gate_3452(G7197,G4083,G4084,G4085,G4086);
nand gate_3453(G986,G984,G985);
nand gate_3454(G989,G987,G988);
nand gate_3455(G1777,G1775,G1776);
nand gate_3456(G1780,G1778,G1779);
not gate_3457(G6259,G6253);
nand gate_3458(G2841,G6253,G6260);
not gate_3459(G7117,G7111);
nand gate_3460(G4077,G7111,G7118);
not gate_3461(G7127,G7121);
nand gate_3462(G4080,G7121,G7128);
nand gate_3463(G6243,G6241,G6242);
not gate_3464(G990,G989);
and gate_3465(G996,G975,G986);
not gate_3466(G1781,G1780);
and gate_3467(G1787,G1766,G1777);
nand gate_3468(G2840,G6256,G6259);
not gate_3469(G6335,G6329);
nand gate_3470(G4076,G7114,G7117);
nand gate_3471(G4079,G7124,G7127);
not gate_3472(G7203,G7197);
and gate_3473(G995,G990,G980);
and gate_3474(G1786,G1781,G1771);
not gate_3475(G6249,G6243);
nand gate_3476(G2838,G6243,G6250);
nand gate_3477(G2842,G2840,G2841);
nand gate_3478(G4078,G4076,G4077);
nand gate_3479(G4081,G4079,G4080);
nand gate_3480(G2837,G6246,G6249);
not gate_3481(G2843,G2842);
not gate_3482(G4082,G4081);
and gate_3483(G4088,G4067,G4078);
or gate_3484(G5170,G995,G996);
or gate_3485(G5740,G1786,G1787);
nand gate_3486(G2839,G2837,G2838);
and gate_3487(G2848,G2843,G2833);
and gate_3488(G4087,G4082,G4072);
nand gate_3489(G1791,G5740,G5743);
nand gate_3490(G1003,G5170,G5173);
not gate_3491(G5174,G5170);
not gate_3492(G5744,G5740);
and gate_3493(G2849,G2828,G2839);
or gate_3494(G7200,G4087,G4088);
nand gate_3495(G1792,G5737,G5744);
nand gate_3496(G1004,G5167,G5174);
or gate_3497(G6332,G2848,G2849);
nand gate_3498(G320,G1791,G1792);
nand gate_3499(G337,G1003,G1004);
nand gate_3500(G4092,G7200,G7203);
not gate_3501(G7204,G7200);
not gate_3502(G321,G320);
not gate_3503(G338,G337);
nand gate_3504(G4093,G7197,G7204);
nand gate_3505(G2855,G6332,G6335);
not gate_3506(G6336,G6332);
nand gate_3507(G369,G4092,G4093);
nand gate_3508(G2856,G6329,G6336);
not gate_3509(G370,G369);
nand gate_3510(G398,G2855,G2856);
not gate_3511(G399,G398);
endmodule
