// Verilog File 
module i8 (pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,po00,po01,po02,po03,po04,po05,
po06,po07,po08,po09,po10,po11,po12,po13,po14,po15,
po16,po17,po18,po19,po20,po21,po22,po23,po24,po25,
po26,po27,po28,po29,po30,po31,po32,po33,po34,po35,
po36,po37,po38,po39,po40,po41,po42,po43,po44,po45,
po46,po47,po48,po49,po50,po51,po52,po53,po54,po55,
po56,po57,po58,po59,po60,po61,po62,po63,po64,po65,
po66,po67,po68,po69,po70,po71,po72,po73,po74,po75,
po76,po77,po78,po79,po80);

input pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18,
po19,po20,po21,po22,po23,po24,po25,po26,po27,po28,
po29,po30,po31,po32,po33,po34,po35,po36,po37,po38,
po39,po40,po41,po42,po43,po44,po45,po46,po47,po48,
po49,po50,po51,po52,po53,po54,po55,po56,po57,po58,
po59,po60,po61,po62,po63,po64,po65,po66,po67,po68,
po69,po70,po71,po72,po73,po74,po75,po76,po77,po78,
po79,po80;

wire n214,n215,n216,n217,n218,n219,n220,n221,n222,
n223,n224,n225,n226,n227,n228,n229,n230,n231,n232,
n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,
n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,
n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,
n263,n264,n266,n267,n268,n269,n270,n271,n272,n273,
n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,
n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,
n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,
n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,
n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,
n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,
n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,
n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,
n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,
n364,n365,n366,n367,n368,n369,n370,n372,n373,n374,
n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,
n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,
n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,
n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,
n415,n416,n417,n419,n420,n421,n422,n423,n424,n425,
n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,
n436,n437,n438,n439,n440,n441,n442,n443,n444,n445,
n446,n447,n448,n449,n450,n451,n452,n453,n454,n455,
n456,n458,n459,n460,n461,n462,n463,n464,n465,n466,
n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,
n477,n478,n479,n480,n481,n483,n484,n485,n486,n487,
n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,
n498,n499,n500,n501,n502,n503,n504,n505,n507,n508,
n509,n510,n511,n512,n513,n514,n515,n516,n517,n518,
n519,n520,n521,n522,n523,n524,n525,n526,n527,n528,
n529,n531,n532,n533,n534,n535,n536,n537,n538,n539,
n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,
n550,n551,n552,n553,n555,n556,n557,n558,n559,n560,
n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,
n571,n572,n573,n574,n575,n576,n577,n579,n580,n581,
n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,
n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,
n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,
n612,n614,n615,n616,n617,n618,n619,n620,n621,n622,
n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,
n633,n634,n635,n636,n637,n638,n639,n641,n642,n643,
n644,n645,n646,n647,n648,n649,n650,n651,n652,n653,
n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,
n664,n665,n666,n667,n669,n670,n671,n672,n673,n674,
n675,n676,n677,n678,n679,n680,n681,n682,n683,n684,
n685,n686,n687,n688,n689,n690,n691,n692,n693,n694,
n695,n696,n697,n698,n699,n700,n701,n702,n703,n704,
n705,n706,n707,n708,n709,n710,n711,n712,n713,n714,
n715,n716,n717,n718,n719,n720,n721,n722,n723,n724,
n726,n727,n728,n729,n730,n731,n732,n733,n734,n735,
n736,n737,n738,n739,n740,n741,n742,n743,n744,n745,
n746,n747,n748,n749,n750,n751,n752,n753,n754,n755,
n756,n757,n758,n759,n760,n761,n762,n763,n764,n765,
n766,n767,n768,n769,n770,n771,n772,n773,n774,n775,
n777,n778,n779,n780,n781,n782,n783,n784,n785,n786,
n787,n788,n789,n790,n791,n792,n793,n794,n795,n796,
n797,n798,n799,n800,n801,n802,n803,n804,n805,n806,
n807,n808,n809,n810,n811,n812,n813,n815,n816,n817,
n818,n819,n820,n821,n822,n823,n824,n825,n826,n827,
n828,n829,n830,n831,n832,n833,n834,n835,n836,n837,
n838,n839,n840,n841,n842,n843,n844,n845,n846,n847,
n848,n849,n850,n851,n853,n854,n855,n856,n857,n858,
n859,n860,n861,n862,n863,n864,n865,n866,n867,n868,
n869,n870,n871,n872,n873,n874,n875,n876,n877,n878,
n879,n880,n881,n882,n883,n884,n885,n886,n887,n888,
n889,n890,n891,n892,n893,n894,n895,n896,n897,n898,
n899,n900,n901,n902,n903,n904,n905,n906,n907,n908,
n909,n911,n912,n913,n914,n915,n916,n917,n918,n919,
n920,n921,n922,n923,n924,n925,n926,n927,n928,n929,
n930,n931,n932,n933,n934,n935,n936,n937,n938,n939,
n940,n941,n942,n943,n944,n945,n946,n947,n949,n950,
n951,n952,n953,n954,n955,n956,n957,n958,n959,n960,
n961,n962,n963,n964,n965,n966,n967,n968,n969,n970,
n971,n972,n973,n974,n975,n976,n977,n978,n979,n980,
n981,n982,n983,n984,n985,n987,n988,n989,n990,n991,
n992,n993,n994,n995,n996,n997,n998,n999,n1000,n1001,
n1002,n1003,n1004,n1005,n1006,n1007,n1008,n1009,n1010,n1011,
n1012,n1013,n1014,n1015,n1016,n1017,n1018,n1019,n1020,n1021,
n1022,n1023,n1025,n1026,n1027,n1028,n1029,n1030,n1031,n1032,
n1033,n1034,n1035,n1036,n1037,n1038,n1039,n1040,n1041,n1042,
n1043,n1044,n1045,n1046,n1047,n1048,n1049,n1050,n1051,n1052,
n1053,n1054,n1055,n1056,n1057,n1058,n1059,n1060,n1061,n1063,
n1064,n1065,n1066,n1067,n1068,n1069,n1070,n1071,n1072,n1073,
n1074,n1075,n1076,n1077,n1078,n1079,n1080,n1081,n1082,n1083,
n1084,n1085,n1086,n1087,n1088,n1089,n1090,n1091,n1092,n1093,
n1094,n1095,n1096,n1097,n1099,n1100,n1101,n1102,n1103,n1104,
n1105,n1106,n1107,n1108,n1109,n1110,n1111,n1112,n1113,n1114,
n1115,n1116,n1117,n1118,n1119,n1120,n1121,n1122,n1123,n1124,
n1125,n1126,n1127,n1128,n1129,n1130,n1131,n1132,n1133,n1135,
n1136,n1137,n1138,n1139,n1140,n1141,n1142,n1143,n1144,n1145,
n1146,n1147,n1148,n1149,n1150,n1151,n1152,n1153,n1154,n1155,
n1156,n1157,n1158,n1159,n1160,n1161,n1162,n1163,n1164,n1165,
n1166,n1167,n1168,n1169,n1171,n1172,n1173,n1174,n1175,n1176,
n1177,n1178,n1179,n1180,n1181,n1182,n1183,n1184,n1185,n1186,
n1187,n1188,n1189,n1190,n1191,n1192,n1193,n1194,n1195,n1196,
n1197,n1198,n1199,n1200,n1201,n1202,n1203,n1204,n1205,n1207,
n1208,n1209,n1210,n1211,n1212,n1213,n1214,n1215,n1216,n1217,
n1218,n1219,n1220,n1221,n1222,n1223,n1224,n1225,n1226,n1227,
n1228,n1229,n1230,n1231,n1232,n1233,n1234,n1235,n1236,n1237,
n1238,n1239,n1240,n1241,n1243,n1244,n1245,n1246,n1247,n1248,
n1249,n1250,n1251,n1252,n1253,n1254,n1255,n1256,n1257,n1258,
n1259,n1260,n1261,n1262,n1263,n1264,n1265,n1266,n1267,n1268,
n1269,n1270,n1271,n1272,n1273,n1274,n1275,n1276,n1277,n1279,
n1280,n1281,n1282,n1283,n1284,n1285,n1286,n1287,n1288,n1289,
n1290,n1291,n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,
n1300,n1301,n1302,n1303,n1304,n1305,n1306,n1307,n1308,n1309,
n1310,n1311,n1312,n1313,n1315,n1316,n1317,n1318,n1319,n1320,
n1321,n1322,n1323,n1324,n1325,n1326,n1327,n1328,n1329,n1330,
n1331,n1332,n1333,n1334,n1335,n1336,n1337,n1338,n1339,n1340,
n1341,n1342,n1343,n1344,n1345,n1346,n1347,n1349,n1350,n1351,
n1352,n1353,n1354,n1355,n1356,n1357,n1358,n1359,n1360,n1361,
n1362,n1363,n1364,n1365,n1366,n1367,n1368,n1369,n1370,n1371,
n1372,n1373,n1374,n1375,n1376,n1377,n1378,n1379,n1380,n1381,
n1383,n1384,n1385,n1386,n1387,n1388,n1389,n1390,n1391,n1392,
n1393,n1394,n1395,n1396,n1397,n1398,n1399,n1400,n1401,n1402,
n1403,n1404,n1405,n1406,n1407,n1408,n1409,n1410,n1411,n1412,
n1413,n1414,n1415,n1417,n1418,n1419,n1420,n1421,n1422,n1423,
n1424,n1425,n1426,n1427,n1428,n1429,n1430,n1431,n1432,n1433,
n1434,n1435,n1436,n1437,n1438,n1439,n1440,n1441,n1442,n1443,
n1444,n1445,n1446,n1447,n1448,n1449,n1451,n1452,n1453,n1454,
n1455,n1456,n1457,n1458,n1459,n1460,n1461,n1462,n1463,n1464,
n1465,n1466,n1467,n1468,n1469,n1470,n1471,n1472,n1473,n1474,
n1475,n1476,n1477,n1478,n1479,n1480,n1481,n1482,n1483,n1484,
n1485,n1486,n1487,n1488,n1489,n1490,n1491,n1492,n1493,n1494,
n1495,n1496,n1497,n1498,n1499,n1500,n1501,n1502,n1503,n1504,
n1505,n1506,n1507,n1508,n1509,n1510,n1511,n1512,n1514,n1515,
n1516,n1517,n1518,n1519,n1520,n1521,n1522,n1523,n1524,n1525,
n1526,n1527,n1528,n1529,n1530,n1531,n1532,n1533,n1534,n1535,
n1536,n1537,n1538,n1539,n1540,n1541,n1542,n1543,n1544,n1545,
n1546,n1547,n1548,n1550,n1551,n1552,n1553,n1554,n1555,n1556,
n1557,n1558,n1559,n1560,n1561,n1562,n1563,n1564,n1565,n1566,
n1567,n1568,n1569,n1570,n1571,n1572,n1573,n1574,n1575,n1576,
n1577,n1578,n1579,n1580,n1581,n1582,n1583,n1584,n1586,n1587,
n1588,n1589,n1590,n1591,n1592,n1593,n1594,n1595,n1596,n1597,
n1598,n1599,n1600,n1601,n1602,n1603,n1604,n1605,n1606,n1607,
n1608,n1609,n1610,n1611,n1612,n1613,n1614,n1615,n1616,n1617,
n1618,n1619,n1620,n1622,n1623,n1624,n1625,n1626,n1627,n1628,
n1629,n1630,n1631,n1632,n1633,n1634,n1635,n1636,n1637,n1638,
n1639,n1640,n1641,n1642,n1643,n1644,n1645,n1646,n1647,n1648,
n1649,n1650,n1651,n1652,n1653,n1654,n1656,n1657,n1658,n1659,
n1660,n1661,n1662,n1663,n1664,n1665,n1666,n1667,n1668,n1669,
n1670,n1671,n1672,n1673,n1674,n1675,n1676,n1677,n1678,n1679,
n1680,n1681,n1682,n1683,n1684,n1685,n1686,n1688,n1689,n1690,
n1691,n1692,n1693,n1694,n1695,n1696,n1697,n1698,n1699,n1700,
n1701,n1702,n1703,n1704,n1705,n1706,n1707,n1708,n1709,n1710,
n1711,n1712,n1713,n1714,n1715,n1716,n1717,n1718,n1720,n1721,
n1722,n1723,n1724,n1725,n1726,n1727,n1728,n1729,n1730,n1731,
n1732,n1733,n1734,n1735,n1736,n1737,n1738,n1739,n1740,n1741,
n1742,n1743,n1744,n1745,n1746,n1747,n1748,n1749,n1750,n1752,
n1753,n1754,n1755,n1756,n1757,n1758,n1759,n1760,n1761,n1762,
n1763,n1764,n1765,n1766,n1767,n1768,n1769,n1770,n1771,n1772,
n1773,n1774,n1775,n1776,n1777,n1778,n1779,n1780,n1781,n1782,
n1784,n1785,n1786,n1787,n1788,n1789,n1790,n1791,n1792,n1793,
n1794,n1795,n1796,n1797,n1798,n1799,n1800,n1801,n1802,n1803,
n1804,n1805,n1806,n1807,n1808,n1809,n1810,n1811,n1812,n1814,
n1815,n1816,n1817,n1818,n1819,n1820,n1821,n1822,n1823,n1824,
n1825,n1826,n1827,n1828,n1829,n1830,n1831,n1832,n1833,n1834,
n1835,n1836,n1837,n1838,n1839,n1840,n1841,n1842,n1844,n1845,
n1846,n1847,n1848,n1849,n1850,n1851,n1852,n1853,n1854,n1855,
n1856,n1857,n1858,n1859,n1860,n1861,n1862,n1863,n1864,n1865,
n1866,n1867,n1868,n1869,n1870,n1871,n1872,n1874,n1875,n1876,
n1877,n1878,n1879,n1880,n1881,n1882,n1883,n1884,n1885,n1886,
n1887,n1888,n1889,n1890,n1891,n1892,n1893,n1894,n1895,n1896,
n1897,n1898,n1899,n1900,n1901,n1902,n1904,n1905,n1906,n1907,
n1908,n1909,n1910,n1911,n1912,n1913,n1914,n1915,n1916,n1917,
n1918,n1919,n1920,n1921,n1922,n1923,n1924,n1925,n1926,n1927,
n1928,n1929,n1930,n1931,n1932,n1934,n1935,n1936,n1937,n1938,
n1939,n1940,n1941,n1942,n1943,n1944,n1945,n1946,n1947,n1948,
n1949,n1950,n1951,n1952,n1953,n1954,n1955,n1956,n1957,n1958,
n1959,n1960,n1961,n1962,n1964,n1965,n1966,n1967,n1968,n1969,
n1970,n1971,n1972,n1973,n1974,n1975,n1976,n1977,n1978,n1979,
n1980,n1981,n1982,n1983,n1984,n1985,n1986,n1987,n1988,n1989,
n1990,n1991,n1992,n1994,n1995,n1996,n1997,n1998,n1999,n2000,
n2001,n2002,n2003,n2004,n2005,n2006,n2007,n2008,n2009,n2010,
n2011,n2012,n2013,n2014,n2015,n2016,n2017,n2018,n2019,n2020,
n2021,n2022,n2023,n2024,n2026,n2027,n2028,n2029,n2030,n2031,
n2032,n2033,n2034,n2035,n2036,n2037,n2038,n2039,n2040,n2041,
n2042,n2043,n2044,n2045,n2046,n2047,n2048,n2049,n2050,n2051,
n2052,n2053,n2054,n2055,n2056,n2058,n2059,n2060,n2061,n2062,
n2063,n2064,n2065,n2066,n2067,n2068,n2069,n2070,n2071,n2072,
n2073,n2074,n2075,n2076,n2077,n2078,n2079,n2080,n2081,n2082,
n2083,n2084,n2085,n2086,n2087,n2088,n2090,n2091,n2092,n2093,
n2094,n2095,n2096,n2097,n2098,n2099,n2100,n2101,n2102,n2103,
n2104,n2105,n2106,n2107,n2108,n2109,n2110,n2111,n2112,n2113,
n2114,n2115,n2116,n2117,n2118,n2119,n2120,n2122,n2123,n2124,
n2125,n2126,n2127,n2128,n2129,n2130,n2131,n2132,n2133,n2134,
n2135,n2136,n2137,n2138,n2139,n2140,n2141,n2142,n2143,n2144,
n2145,n2146,n2147,n2148,n2149,n2150,n2151,n2152,n2153,n2154,
n2156,n2157,n2158,n2159,n2160,n2161,n2162,n2163,n2164,n2165,
n2166,n2167,n2168,n2169,n2170,n2171,n2172,n2173,n2174,n2175,
n2176,n2177,n2178,n2179,n2180,n2181,n2182,n2183,n2184,n2185,
n2186,n2188,n2189,n2190,n2191,n2192,n2193,n2194,n2195,n2196,
n2197,n2198,n2199,n2200,n2201,n2202,n2203,n2204,n2205,n2206,
n2207,n2208,n2209,n2210,n2211,n2212,n2213,n2214,n2215,n2216,
n2217,n2218,n2220,n2221,n2222,n2223,n2224,n2225,n2226,n2227,
n2228,n2229,n2230,n2231,n2232,n2233,n2234,n2235,n2236,n2237,
n2238,n2239,n2240,n2241,n2242,n2243,n2244,n2245,n2246,n2247,
n2248,n2249,n2250,n2251,n2253,n2254,n2255,n2256,n2257,n2258,
n2259,n2260,n2261,n2262,n2263,n2264,n2265,n2266,n2267,n2268,
n2269,n2270,n2271,n2272,n2273,n2274,n2275,n2276,n2277,n2278,
n2279,n2280,n2281,n2282,n2283,n2284,n2286,n2287,n2288,n2289,
n2290,n2291,n2292,n2293,n2294,n2295,n2296,n2297,n2298,n2299,
n2300,n2301,n2302,n2303,n2304,n2305,n2306,n2307,n2308,n2309,
n2310,n2311,n2312,n2313,n2314,n2315,n2316,n2318,n2319,n2320,
n2321,n2322,n2323,n2324,n2325,n2326,n2327,n2328,n2329,n2330,
n2331,n2332,n2333,n2334,n2335,n2336,n2337,n2338,n2339,n2340,
n2341,n2342,n2343,n2344,n2345,n2346,n2347,n2348,n2350,n2351,
n2352,n2353,n2354,n2355,n2356,n2357,n2358,n2359,n2360,n2361,
n2362,n2363,n2364,n2365,n2366,n2367,n2368,n2369,n2370,n2371,
n2372,n2373,n2374,n2375,n2376,n2377,n2378,n2379,n2380,n2382,
n2383,n2384,n2385,n2386,n2387,n2388,n2389,n2390,n2391,n2392,
n2393,n2394,n2395,n2396,n2397,n2398,n2399,n2400,n2401,n2402,
n2403,n2404,n2405,n2406,n2407,n2408,n2409,n2410,n2412,n2413,
n2414,n2415,n2416,n2417,n2418,n2419,n2420,n2421,n2422,n2423,
n2424,n2425,n2426,n2427,n2428,n2429,n2430,n2431,n2432,n2433,
n2434,n2435,n2436,n2437,n2438,n2439,n2440,n2441,n2443,n2444,
n2445,n2446,n2447,n2448,n2449,n2450,n2451,n2452,n2453,n2454,
n2455,n2456,n2457,n2458,n2459,n2460,n2461,n2462,n2463,n2464,
n2465,n2466,n2467,n2468,n2469,n2470,n2471,n2472,n2474,n2475,
n2476,n2477,n2478,n2479,n2480,n2481,n2482,n2483,n2484,n2485,
n2486,n2487,n2488,n2489,n2490,n2491,n2492,n2493,n2494,n2495,
n2496,n2497,n2498,n2499,n2500,n2501,n2502,n2503,n2505,n2506,
n2507,n2508,n2509,n2510,n2511,n2512,n2513,n2514,n2515,n2516,
n2517,n2518,n2519,n2520,n2521,n2522,n2523,n2524,n2525,n2526,
n2527,n2529,n2530,n2531,n2532,n2533,n2534,n2535,n2537,n2538,
n2539,n2540,n2541,n2542,n2543,n2545,n2546,n2547,n2548,n2549,
n2550,n2551,n2553,n2554,n2555,n2556,n2557,n2558,n2559,n2561,
n2562,n2563,n2564,n2565,n2566,n2567,n2569,n2570,n2571,n2572,
n2573,n2574,n2575,n2577,n2578,n2579,n2580,n2581,n2582,n2583,
n2585,n2586,n2587,n2588,n2589,n2590,n2591,n2593,n2594,n2595,
n2596,n2597,n2598,n2599,n2601,n2602,n2603,n2604,n2605,n2606,
n2607,n2609,n2610,n2611,n2612,n2613,n2614,n2615,n2617,n2618,
n2619,n2620,n2621,n2622,n2623,n2625,n2626,n2627,n2628,n2629,
n2630,n2631,n2633,n2634,n2635,n2636,n2637,n2638,n2639,n2641,
n2642,n2643,n2644,n2645,n2646,n2647,n2648,n2649,n2650,n2651,
n2652,n2653,n2654,n2655,n2656,n2657,n2658,n2659,n2660,n2661,
n2662,n2663,n2664,n2666,n2667,n2668,n2669,n2670,n2671,n2672,
n2673,n2674,n2675,n2676;
not gate_0(n214,pi000);
not gate_1(n215,pi001);
not gate_2(n216,pi002);
not gate_3(n217,pi003);
not gate_4(n218,pi004);
not gate_5(n219,pi005);
not gate_6(n220,pi006);
not gate_7(n221,pi007);
not gate_8(n222,pi008);
not gate_9(n223,pi095);
not gate_10(n224,pi130);
not gate_11(n225,pi131);
not gate_12(n226,pi132);
and gate_13(n227,n219,n223);
and gate_14(n228,n221,n227);
not gate_15(n229,n228);
and gate_16(n230,n216,n227);
and gate_17(n231,pi007,n230);
not gate_18(n232,n231);
and gate_19(n233,pi089,n232);
and gate_20(n234,n228,n233);
not gate_21(n235,n234);
and gate_22(n236,n215,n219);
and gate_23(n237,n223,n236);
and gate_24(n238,pi007,n237);
not gate_25(n239,n238);
and gate_26(n240,n232,n239);
not gate_27(n241,n240);
and gate_28(n242,pi088,n241);
not gate_29(n243,n242);
and gate_30(n244,n235,n243);
and gate_31(n245,n219,pi095);
not gate_32(n246,n245);
and gate_33(n247,n219,n229);
and gate_34(n248,n239,n247);
and gate_35(n249,n232,n248);
and gate_36(n250,n246,n249);
not gate_37(n251,n250);
and gate_38(n252,pi090,n229);
and gate_39(n253,n239,n252);
and gate_40(n254,n232,n253);
and gate_41(n255,n245,n254);
not gate_42(n256,n255);
and gate_43(n257,pi087,n246);
and gate_44(n258,n232,n257);
and gate_45(n259,n239,n258);
and gate_46(n260,pi005,n259);
not gate_47(n261,n260);
and gate_48(n262,n256,n261);
and gate_49(n263,n251,n262);
and gate_50(n264,n244,n263);
not gate_51(po00,n264);
and gate_52(n266,n221,n230);
not gate_53(n267,n266);
and gate_54(n268,pi008,n227);
not gate_55(n269,n268);
and gate_56(n270,n222,n223);
and gate_57(n271,pi007,n270);
not gate_58(n272,n271);
and gate_59(n273,pi001,n223);
and gate_60(n274,pi002,n273);
and gate_61(n275,n222,n274);
and gate_62(n276,n224,n275);
not gate_63(n277,n276);
and gate_64(n278,n221,n237);
not gate_65(n279,n278);
and gate_66(n280,n219,n279);
and gate_67(n281,pi092,n280);
and gate_68(n282,n277,n281);
and gate_69(n283,n272,n282);
and gate_70(n284,n269,n283);
and gate_71(n285,n266,n284);
not gate_72(n286,n285);
and gate_73(n287,pi094,n267);
and gate_74(n288,n269,n287);
and gate_75(n289,n272,n288);
and gate_76(n290,n277,n289);
and gate_77(n291,n280,n290);
and gate_78(n292,n245,n291);
not gate_79(n293,n292);
and gate_80(n294,pi092,n269);
and gate_81(n295,n272,n294);
and gate_82(n296,n277,n295);
and gate_83(n297,n278,n296);
not gate_84(n298,n297);
and gate_85(n299,n293,n298);
and gate_86(n300,n286,n299);
and gate_87(n301,pi000,pi001);
and gate_88(n302,pi002,n301);
not gate_89(n303,n302);
and gate_90(n304,n219,n303);
not gate_91(n305,n304);
and gate_92(n306,pi038,n305);
not gate_93(n307,n306);
and gate_94(n308,n218,n219);
and gate_95(n309,n215,n308);
and gate_96(n310,pi003,n309);
and gate_97(n311,pi002,n310);
and gate_98(n312,n220,n311);
not gate_99(n313,n312);
and gate_100(n314,pi002,n219);
and gate_101(n315,n215,n314);
and gate_102(n316,pi008,n315);
not gate_103(n317,n316);
and gate_104(n318,pi001,n219);
and gate_105(n319,pi002,n318);
not gate_106(n320,n319);
and gate_107(n321,n214,n319);
not gate_108(n322,n321);
and gate_109(n323,n317,n322);
and gate_110(n324,n313,n323);
not gate_111(n325,n324);
and gate_112(n326,n216,n309);
and gate_113(n327,n220,n326);
not gate_114(n328,n327);
and gate_115(n329,n216,pi007);
and gate_116(n330,n236,n329);
not gate_117(n331,n330);
and gate_118(n332,n328,n331);
not gate_119(n333,n332);
and gate_120(n334,pi008,n318);
not gate_121(n335,n334);
and gate_122(n336,pi001,n308);
and gate_123(n337,n216,n336);
and gate_124(n338,n220,n337);
not gate_125(n339,n338);
and gate_126(n340,n335,n339);
and gate_127(n341,n217,n219);
and gate_128(n342,pi004,n221);
not gate_129(n343,n342);
and gate_130(n344,n341,n343);
not gate_131(n345,n344);
and gate_132(n346,n340,n345);
not gate_133(n347,n346);
and gate_134(n348,n332,n346);
and gate_135(n349,n304,n348);
and gate_136(n350,n324,n349);
not gate_137(n351,n350);
and gate_138(n352,n307,n351);
and gate_139(n353,pi050,n346);
and gate_140(n354,n304,n353);
and gate_141(n355,n325,n354);
not gate_142(n356,n355);
and gate_143(n357,pi065,n324);
and gate_144(n358,n304,n357);
and gate_145(n359,n346,n358);
and gate_146(n360,n333,n359);
not gate_147(n361,n360);
and gate_148(n362,n356,n361);
and gate_149(n363,n352,n362);
not gate_150(n364,n363);
and gate_151(n365,n219,n277);
and gate_152(n366,n272,n365);
not gate_153(n367,n366);
and gate_154(n368,n364,n367);
not gate_155(n369,n368);
and gate_156(n370,n300,n369);
not gate_157(po01,n370);
and gate_158(n372,pi039,n305);
not gate_159(n373,n372);
and gate_160(n374,n351,n373);
and gate_161(n375,pi051,n346);
and gate_162(n376,n304,n375);
and gate_163(n377,n325,n376);
not gate_164(n378,n377);
and gate_165(n379,pi066,n324);
and gate_166(n380,n304,n379);
and gate_167(n381,n346,n380);
and gate_168(n382,n333,n381);
not gate_169(n383,n382);
and gate_170(n384,n378,n383);
and gate_171(n385,n374,n384);
not gate_172(n386,n385);
and gate_173(n387,n272,n386);
and gate_174(n388,n277,n387);
and gate_175(n389,pi005,n388);
not gate_176(n390,n389);
and gate_177(n391,pi091,n366);
and gate_178(n392,n268,n391);
not gate_179(n393,n392);
and gate_180(n394,n390,n393);
and gate_181(n395,n272,n277);
not gate_182(n396,n395);
and gate_183(n397,n386,n396);
not gate_184(n398,n397);
and gate_185(n399,n394,n398);
and gate_186(n400,pi093,n269);
and gate_187(n401,n366,n400);
and gate_188(n402,n278,n401);
not gate_189(n403,n402);
and gate_190(n404,pi093,n280);
and gate_191(n405,n277,n404);
and gate_192(n406,n272,n405);
and gate_193(n407,n269,n406);
and gate_194(n408,n266,n407);
not gate_195(n409,n408);
and gate_196(n410,n403,n409);
and gate_197(n411,pi096,n267);
and gate_198(n412,n269,n411);
and gate_199(n413,n366,n412);
and gate_200(n414,n245,n413);
not gate_201(n415,n414);
and gate_202(n416,n410,n415);
and gate_203(n417,n399,n416);
not gate_204(po02,n417);
and gate_205(n419,n220,n223);
and gate_206(n420,n224,n419);
not gate_207(n421,n420);
and gate_208(n422,pi044,n346);
and gate_209(n423,n304,n422);
and gate_210(n424,n325,n423);
not gate_211(n425,n424);
and gate_212(n426,pi032,n305);
not gate_213(n427,n426);
and gate_214(n428,pi040,n347);
and gate_215(n429,n304,n428);
not gate_216(n430,n429);
and gate_217(n431,n427,n430);
and gate_218(n432,n425,n431);
and gate_219(n433,pi059,n324);
and gate_220(n434,n304,n433);
and gate_221(n435,n346,n434);
and gate_222(n436,n333,n435);
not gate_223(n437,n436);
and gate_224(n438,n351,n437);
and gate_225(n439,n432,n438);
not gate_226(n440,n439);
and gate_227(n441,pi007,n223);
not gate_228(n442,n441);
and gate_229(n443,n440,n442);
and gate_230(n444,n421,n443);
and gate_231(n445,pi005,n444);
not gate_232(n446,n445);
and gate_233(n447,n219,pi097);
and gate_234(n448,n421,n447);
and gate_235(n449,n245,n448);
not gate_236(n450,n449);
and gate_237(n451,n446,n450);
and gate_238(n452,n421,n442);
not gate_239(n453,n452);
and gate_240(n454,n440,n453);
not gate_241(n455,n454);
and gate_242(n456,n451,n455);
not gate_243(po03,n456);
and gate_244(n458,n219,pi098);
and gate_245(n459,n452,n458);
and gate_246(n460,n245,n459);
not gate_247(n461,n460);
and gate_248(n462,pi033,n305);
not gate_249(n463,n462);
and gate_250(n464,n351,n463);
and gate_251(n465,pi045,n346);
and gate_252(n466,n304,n465);
and gate_253(n467,n325,n466);
not gate_254(n468,n467);
and gate_255(n469,pi060,n324);
and gate_256(n470,n304,n469);
and gate_257(n471,n346,n470);
and gate_258(n472,n333,n471);
not gate_259(n473,n472);
and gate_260(n474,n468,n473);
and gate_261(n475,n464,n474);
not gate_262(n476,n475);
and gate_263(n477,n219,n452);
not gate_264(n478,n477);
and gate_265(n479,n476,n478);
not gate_266(n480,n479);
and gate_267(n481,n461,n480);
not gate_268(po04,n481);
and gate_269(n483,n219,pi099);
and gate_270(n484,pi095,n483);
not gate_271(n485,n484);
and gate_272(n486,n477,n484);
not gate_273(n487,n486);
and gate_274(n488,pi034,n305);
not gate_275(n489,n488);
and gate_276(n490,n351,n489);
and gate_277(n491,pi046,n346);
and gate_278(n492,n304,n491);
and gate_279(n493,n325,n492);
not gate_280(n494,n493);
and gate_281(n495,pi061,n324);
and gate_282(n496,n304,n495);
and gate_283(n497,n346,n496);
and gate_284(n498,n333,n497);
not gate_285(n499,n498);
and gate_286(n500,n494,n499);
and gate_287(n501,n490,n500);
not gate_288(n502,n501);
and gate_289(n503,n478,n502);
not gate_290(n504,n503);
and gate_291(n505,n487,n504);
not gate_292(po05,n505);
and gate_293(n507,n219,pi100);
and gate_294(n508,pi095,n507);
not gate_295(n509,n508);
and gate_296(n510,n477,n508);
not gate_297(n511,n510);
and gate_298(n512,pi035,n305);
not gate_299(n513,n512);
and gate_300(n514,n351,n513);
and gate_301(n515,pi047,n346);
and gate_302(n516,n304,n515);
and gate_303(n517,n325,n516);
not gate_304(n518,n517);
and gate_305(n519,pi062,n324);
and gate_306(n520,n304,n519);
and gate_307(n521,n346,n520);
and gate_308(n522,n333,n521);
not gate_309(n523,n522);
and gate_310(n524,n518,n523);
and gate_311(n525,n514,n524);
not gate_312(n526,n525);
and gate_313(n527,n478,n526);
not gate_314(n528,n527);
and gate_315(n529,n511,n528);
not gate_316(po06,n529);
and gate_317(n531,n219,pi101);
and gate_318(n532,pi095,n531);
not gate_319(n533,n532);
and gate_320(n534,n477,n532);
not gate_321(n535,n534);
and gate_322(n536,pi036,n305);
not gate_323(n537,n536);
and gate_324(n538,n351,n537);
and gate_325(n539,pi048,n346);
and gate_326(n540,n304,n539);
and gate_327(n541,n325,n540);
not gate_328(n542,n541);
and gate_329(n543,pi063,n324);
and gate_330(n544,n304,n543);
and gate_331(n545,n346,n544);
and gate_332(n546,n333,n545);
not gate_333(n547,n546);
and gate_334(n548,n542,n547);
and gate_335(n549,n538,n548);
not gate_336(n550,n549);
and gate_337(n551,n478,n550);
not gate_338(n552,n551);
and gate_339(n553,n535,n552);
not gate_340(po07,n553);
and gate_341(n555,n219,pi102);
and gate_342(n556,pi095,n555);
not gate_343(n557,n556);
and gate_344(n558,n477,n556);
not gate_345(n559,n558);
and gate_346(n560,pi037,n305);
not gate_347(n561,n560);
and gate_348(n562,n351,n561);
and gate_349(n563,pi049,n346);
and gate_350(n564,n304,n563);
and gate_351(n565,n325,n564);
not gate_352(n566,n565);
and gate_353(n567,pi064,n324);
and gate_354(n568,n304,n567);
and gate_355(n569,n346,n568);
and gate_356(n570,n333,n569);
not gate_357(n571,n570);
and gate_358(n572,n566,n571);
and gate_359(n573,n562,n572);
not gate_360(n574,n573);
and gate_361(n575,n478,n574);
not gate_362(n576,n575);
and gate_363(n577,n559,n576);
not gate_364(po08,n577);
and gate_365(n579,pi043,n346);
and gate_366(n580,n304,n579);
and gate_367(n581,n325,n580);
not gate_368(n582,n581);
and gate_369(n583,pi031,n305);
not gate_370(n584,n583);
and gate_371(n585,pi039,n347);
and gate_372(n586,n304,n585);
not gate_373(n587,n586);
and gate_374(n588,n584,n587);
and gate_375(n589,n582,n588);
and gate_376(n590,pi058,n324);
and gate_377(n591,n304,n590);
and gate_378(n592,n346,n591);
and gate_379(n593,n333,n592);
not gate_380(n594,n593);
and gate_381(n595,n351,n594);
and gate_382(n596,n589,n595);
not gate_383(n597,n596);
and gate_384(n598,n223,n224);
not gate_385(n599,n598);
and gate_386(n600,n442,n599);
not gate_387(n601,n600);
and gate_388(n602,n597,n601);
not gate_389(n603,n602);
and gate_390(n604,n442,n597);
and gate_391(n605,n599,n604);
and gate_392(n606,pi005,n605);
not gate_393(n607,n606);
and gate_394(n608,n219,pi103);
and gate_395(n609,n245,n608);
not gate_396(n610,n609);
and gate_397(n611,n607,n610);
and gate_398(n612,n603,n611);
not gate_399(po09,n612);
and gate_400(n614,n219,pi104);
and gate_401(n615,pi095,n614);
and gate_402(n616,n477,n615);
not gate_403(n617,n616);
and gate_404(n618,pi041,n346);
and gate_405(n619,n304,n618);
and gate_406(n620,n325,n619);
not gate_407(n621,n620);
and gate_408(n622,pi029,n305);
not gate_409(n623,n622);
and gate_410(n624,pi037,n347);
and gate_411(n625,n304,n624);
not gate_412(n626,n625);
and gate_413(n627,n623,n626);
and gate_414(n628,n621,n627);
and gate_415(n629,pi056,n324);
and gate_416(n630,n304,n629);
and gate_417(n631,n346,n630);
and gate_418(n632,n333,n631);
not gate_419(n633,n632);
and gate_420(n634,n351,n633);
and gate_421(n635,n628,n634);
not gate_422(n636,n635);
and gate_423(n637,n478,n636);
not gate_424(n638,n637);
and gate_425(n639,n617,n638);
not gate_426(po10,n639);
and gate_427(n641,n219,pi105);
and gate_428(n642,pi095,n641);
not gate_429(n643,n642);
and gate_430(n644,n477,n642);
not gate_431(n645,n644);
and gate_432(n646,pi042,n346);
and gate_433(n647,n304,n646);
and gate_434(n648,n325,n647);
not gate_435(n649,n648);
and gate_436(n650,pi030,n305);
not gate_437(n651,n650);
and gate_438(n652,pi038,n347);
and gate_439(n653,n304,n652);
not gate_440(n654,n653);
and gate_441(n655,n651,n654);
and gate_442(n656,n649,n655);
and gate_443(n657,pi057,n324);
and gate_444(n658,n304,n657);
and gate_445(n659,n346,n658);
and gate_446(n660,n333,n659);
not gate_447(n661,n660);
and gate_448(n662,n351,n661);
and gate_449(n663,n656,n662);
not gate_450(n664,n663);
and gate_451(n665,n478,n664);
not gate_452(n666,n665);
and gate_453(n667,n645,n666);
not gate_454(po11,n667);
and gate_455(n669,pi039,n346);
and gate_456(n670,n304,n669);
and gate_457(n671,n325,n670);
not gate_458(n672,n671);
and gate_459(n673,pi028,n305);
not gate_460(n674,n673);
and gate_461(n675,pi036,n347);
and gate_462(n676,n304,n675);
not gate_463(n677,n676);
and gate_464(n678,n674,n677);
and gate_465(n679,n672,n678);
and gate_466(n680,pi055,n324);
and gate_467(n681,n304,n680);
and gate_468(n682,n346,n681);
and gate_469(n683,n333,n682);
not gate_470(n684,n683);
and gate_471(n685,n351,n684);
and gate_472(n686,n679,n685);
not gate_473(n687,n686);
and gate_474(n688,n215,n223);
and gate_475(n689,n224,n688);
not gate_476(n690,n689);
and gate_477(n691,n216,n420);
not gate_478(n692,n691);
and gate_479(n693,n690,n692);
and gate_480(n694,pi000,n598);
not gate_481(n695,n694);
and gate_482(n696,n442,n695);
and gate_483(n697,n693,n696);
not gate_484(n698,n697);
and gate_485(n699,n687,n698);
not gate_486(n700,n699);
and gate_487(n701,n687,n692);
and gate_488(n702,n690,n701);
and gate_489(n703,n695,n702);
and gate_490(n704,n442,n703);
and gate_491(n705,pi005,n704);
not gate_492(n706,n705);
and gate_493(n707,n219,pi106);
and gate_494(n708,n695,n707);
and gate_495(n709,n690,n708);
and gate_496(n710,n692,n709);
and gate_497(n711,n245,n710);
not gate_498(n712,n711);
and gate_499(n713,n706,n712);
and gate_500(n714,pi086,n246);
and gate_501(n715,n442,n714);
and gate_502(n716,n692,n715);
and gate_503(n717,n690,n716);
and gate_504(n718,n695,n717);
and gate_505(n719,n228,n718);
and gate_506(n720,n224,n719);
and gate_507(n721,n321,n720);
not gate_508(n722,n721);
and gate_509(n723,n713,n722);
and gate_510(n724,n700,n723);
not gate_511(po12,n724);
and gate_512(n726,pi036,n346);
and gate_513(n727,n304,n726);
and gate_514(n728,n325,n727);
not gate_515(n729,n728);
and gate_516(n730,pi025,n305);
not gate_517(n731,n730);
and gate_518(n732,pi033,n347);
and gate_519(n733,n304,n732);
not gate_520(n734,n733);
and gate_521(n735,n731,n734);
and gate_522(n736,n729,n735);
and gate_523(n737,pi052,n324);
and gate_524(n738,n304,n737);
and gate_525(n739,n346,n738);
and gate_526(n740,n333,n739);
not gate_527(n741,n740);
and gate_528(n742,n351,n741);
and gate_529(n743,n736,n742);
not gate_530(n744,n743);
and gate_531(n745,n220,n688);
and gate_532(n746,n224,n745);
not gate_533(n747,n746);
and gate_534(n748,n692,n747);
and gate_535(n749,n696,n748);
not gate_536(n750,n749);
and gate_537(n751,n744,n750);
not gate_538(n752,n751);
and gate_539(n753,n692,n744);
and gate_540(n754,n747,n753);
and gate_541(n755,n696,n754);
and gate_542(n756,pi005,n755);
not gate_543(n757,n756);
and gate_544(n758,n219,pi107);
and gate_545(n759,n695,n758);
and gate_546(n760,n747,n759);
and gate_547(n761,n692,n760);
and gate_548(n762,n245,n761);
not gate_549(n763,n762);
and gate_550(n764,n757,n763);
and gate_551(n765,pi083,n246);
and gate_552(n766,n442,n765);
and gate_553(n767,n692,n766);
and gate_554(n768,n747,n767);
and gate_555(n769,n695,n768);
and gate_556(n770,n228,n769);
and gate_557(n771,n224,n770);
and gate_558(n772,n321,n771);
not gate_559(n773,n772);
and gate_560(n774,n764,n773);
and gate_561(n775,n752,n774);
not gate_562(po13,n775);
and gate_563(n777,pi037,n346);
and gate_564(n778,n304,n777);
and gate_565(n779,n325,n778);
not gate_566(n780,n779);
and gate_567(n781,pi026,n305);
not gate_568(n782,n781);
and gate_569(n783,pi034,n347);
and gate_570(n784,n304,n783);
not gate_571(n785,n784);
and gate_572(n786,n782,n785);
and gate_573(n787,n780,n786);
and gate_574(n788,pi053,n324);
and gate_575(n789,n304,n788);
and gate_576(n790,n346,n789);
and gate_577(n791,n333,n790);
not gate_578(n792,n791);
and gate_579(n793,n351,n792);
and gate_580(n794,n787,n793);
not gate_581(n795,n794);
and gate_582(n796,n750,n795);
not gate_583(n797,n796);
and gate_584(n798,n748,n795);
and gate_585(n799,n696,n798);
and gate_586(n800,pi005,n799);
not gate_587(n801,n800);
and gate_588(n802,n219,pi108);
and gate_589(n803,n749,n802);
and gate_590(n804,n245,n803);
not gate_591(n805,n804);
and gate_592(n806,n801,n805);
and gate_593(n807,pi084,n749);
and gate_594(n808,n228,n807);
and gate_595(n809,n224,n808);
and gate_596(n810,n321,n809);
not gate_597(n811,n810);
and gate_598(n812,n806,n811);
and gate_599(n813,n797,n812);
not gate_600(po14,n813);
and gate_601(n815,pi038,n346);
and gate_602(n816,n304,n815);
and gate_603(n817,n325,n816);
not gate_604(n818,n817);
and gate_605(n819,pi027,n305);
not gate_606(n820,n819);
and gate_607(n821,pi035,n347);
and gate_608(n822,n304,n821);
not gate_609(n823,n822);
and gate_610(n824,n820,n823);
and gate_611(n825,n818,n824);
and gate_612(n826,pi054,n324);
and gate_613(n827,n304,n826);
and gate_614(n828,n346,n827);
and gate_615(n829,n333,n828);
not gate_616(n830,n829);
and gate_617(n831,n351,n830);
and gate_618(n832,n825,n831);
not gate_619(n833,n832);
and gate_620(n834,n750,n833);
not gate_621(n835,n834);
and gate_622(n836,n748,n833);
and gate_623(n837,n696,n836);
and gate_624(n838,pi005,n837);
not gate_625(n839,n838);
and gate_626(n840,n219,pi109);
and gate_627(n841,n749,n840);
and gate_628(n842,n245,n841);
not gate_629(n843,n842);
and gate_630(n844,n839,n843);
and gate_631(n845,pi085,n749);
and gate_632(n846,n228,n845);
and gate_633(n847,n224,n846);
and gate_634(n848,n321,n847);
not gate_635(n849,n848);
and gate_636(n850,n844,n849);
and gate_637(n851,n835,n850);
not gate_638(po15,n851);
and gate_639(n853,n216,n688);
and gate_640(n854,n224,n853);
not gate_641(n855,n854);
and gate_642(n856,pi035,n346);
and gate_643(n857,n304,n856);
and gate_644(n858,n325,n857);
not gate_645(n859,n858);
and gate_646(n860,pi024,n305);
not gate_647(n861,n860);
and gate_648(n862,pi032,n347);
and gate_649(n863,n304,n862);
not gate_650(n864,n863);
and gate_651(n865,n861,n864);
and gate_652(n866,n859,n865);
and gate_653(n867,n324,n670);
and gate_654(n868,n333,n867);
not gate_655(n869,n868);
and gate_656(n870,n351,n869);
and gate_657(n871,n866,n870);
not gate_658(n872,n871);
and gate_659(n873,n747,n872);
and gate_660(n874,n855,n873);
and gate_661(n875,n692,n874);
and gate_662(n876,n695,n875);
and gate_663(n877,n441,n876);
not gate_664(n878,n877);
and gate_665(n879,n442,n872);
and gate_666(n880,n855,n879);
and gate_667(n881,n748,n880);
and gate_668(n882,n695,n881);
and gate_669(n883,pi005,n882);
not gate_670(n884,n883);
and gate_671(n885,n878,n884);
and gate_672(n886,n219,pi110);
and gate_673(n887,n695,n886);
and gate_674(n888,n855,n887);
and gate_675(n889,n748,n888);
and gate_676(n890,n245,n889);
not gate_677(n891,n890);
and gate_678(n892,pi082,n246);
and gate_679(n893,n442,n892);
and gate_680(n894,n855,n893);
and gate_681(n895,n748,n894);
and gate_682(n896,n695,n895);
and gate_683(n897,n228,n896);
and gate_684(n898,n224,n897);
and gate_685(n899,n321,n898);
not gate_686(n900,n899);
and gate_687(n901,n891,n900);
and gate_688(n902,n885,n901);
and gate_689(n903,n747,n855);
and gate_690(n904,n692,n695);
and gate_691(n905,n903,n904);
not gate_692(n906,n905);
and gate_693(n907,n872,n906);
not gate_694(n908,n907);
and gate_695(n909,n902,n908);
not gate_696(po16,n909);
and gate_697(n911,pi020,n346);
and gate_698(n912,n304,n911);
and gate_699(n913,n325,n912);
not gate_700(n914,n913);
and gate_701(n915,pi009,n305);
not gate_702(n916,n915);
and gate_703(n917,pi017,n347);
and gate_704(n918,n304,n917);
not gate_705(n919,n918);
and gate_706(n920,n916,n919);
and gate_707(n921,n914,n920);
and gate_708(n922,pi024,n346);
and gate_709(n923,n304,n922);
and gate_710(n924,n324,n923);
and gate_711(n925,n333,n924);
not gate_712(n926,n925);
and gate_713(n927,n351,n926);
and gate_714(n928,n921,n927);
not gate_715(n929,n928);
and gate_716(n930,n750,n929);
not gate_717(n931,n930);
and gate_718(n932,n748,n929);
and gate_719(n933,n696,n932);
and gate_720(n934,pi005,n933);
not gate_721(n935,n934);
and gate_722(n936,n219,pi111);
and gate_723(n937,n749,n936);
and gate_724(n938,n245,n937);
not gate_725(n939,n938);
and gate_726(n940,n935,n939);
and gate_727(n941,pi067,n749);
and gate_728(n942,n228,n941);
and gate_729(n943,n224,n942);
and gate_730(n944,n321,n943);
not gate_731(n945,n944);
and gate_732(n946,n940,n945);
and gate_733(n947,n931,n946);
not gate_734(po17,n947);
and gate_735(n949,pi021,n346);
and gate_736(n950,n304,n949);
and gate_737(n951,n325,n950);
not gate_738(n952,n951);
and gate_739(n953,pi010,n305);
not gate_740(n954,n953);
and gate_741(n955,pi018,n347);
and gate_742(n956,n304,n955);
not gate_743(n957,n956);
and gate_744(n958,n954,n957);
and gate_745(n959,n952,n958);
and gate_746(n960,pi025,n346);
and gate_747(n961,n304,n960);
and gate_748(n962,n324,n961);
and gate_749(n963,n333,n962);
not gate_750(n964,n963);
and gate_751(n965,n351,n964);
and gate_752(n966,n959,n965);
not gate_753(n967,n966);
and gate_754(n968,n750,n967);
not gate_755(n969,n968);
and gate_756(n970,n748,n967);
and gate_757(n971,n696,n970);
and gate_758(n972,pi005,n971);
not gate_759(n973,n972);
and gate_760(n974,n219,pi112);
and gate_761(n975,n749,n974);
and gate_762(n976,n245,n975);
not gate_763(n977,n976);
and gate_764(n978,n973,n977);
and gate_765(n979,pi068,n749);
and gate_766(n980,n228,n979);
and gate_767(n981,n224,n980);
and gate_768(n982,n321,n981);
not gate_769(n983,n982);
and gate_770(n984,n978,n983);
and gate_771(n985,n969,n984);
not gate_772(po18,n985);
and gate_773(n987,pi022,n346);
and gate_774(n988,n304,n987);
and gate_775(n989,n325,n988);
not gate_776(n990,n989);
and gate_777(n991,pi011,n305);
not gate_778(n992,n991);
and gate_779(n993,pi019,n347);
and gate_780(n994,n304,n993);
not gate_781(n995,n994);
and gate_782(n996,n992,n995);
and gate_783(n997,n990,n996);
and gate_784(n998,pi026,n346);
and gate_785(n999,n304,n998);
and gate_786(n1000,n324,n999);
and gate_787(n1001,n333,n1000);
not gate_788(n1002,n1001);
and gate_789(n1003,n351,n1002);
and gate_790(n1004,n997,n1003);
not gate_791(n1005,n1004);
and gate_792(n1006,n750,n1005);
not gate_793(n1007,n1006);
and gate_794(n1008,n748,n1005);
and gate_795(n1009,n696,n1008);
and gate_796(n1010,pi005,n1009);
not gate_797(n1011,n1010);
and gate_798(n1012,n219,pi113);
and gate_799(n1013,n749,n1012);
and gate_800(n1014,n245,n1013);
not gate_801(n1015,n1014);
and gate_802(n1016,n1011,n1015);
and gate_803(n1017,pi069,n749);
and gate_804(n1018,n228,n1017);
and gate_805(n1019,n224,n1018);
and gate_806(n1020,n321,n1019);
not gate_807(n1021,n1020);
and gate_808(n1022,n1016,n1021);
and gate_809(n1023,n1007,n1022);
not gate_810(po19,n1023);
and gate_811(n1025,pi023,n346);
and gate_812(n1026,n304,n1025);
and gate_813(n1027,n325,n1026);
not gate_814(n1028,n1027);
and gate_815(n1029,pi012,n305);
not gate_816(n1030,n1029);
and gate_817(n1031,pi020,n347);
and gate_818(n1032,n304,n1031);
not gate_819(n1033,n1032);
and gate_820(n1034,n1030,n1033);
and gate_821(n1035,n1028,n1034);
and gate_822(n1036,pi027,n346);
and gate_823(n1037,n304,n1036);
and gate_824(n1038,n324,n1037);
and gate_825(n1039,n333,n1038);
not gate_826(n1040,n1039);
and gate_827(n1041,n351,n1040);
and gate_828(n1042,n1035,n1041);
not gate_829(n1043,n1042);
and gate_830(n1044,n750,n1043);
not gate_831(n1045,n1044);
and gate_832(n1046,n748,n1043);
and gate_833(n1047,n696,n1046);
and gate_834(n1048,pi005,n1047);
not gate_835(n1049,n1048);
and gate_836(n1050,n219,pi114);
and gate_837(n1051,n749,n1050);
and gate_838(n1052,n245,n1051);
not gate_839(n1053,n1052);
and gate_840(n1054,n1049,n1053);
and gate_841(n1055,pi070,n749);
and gate_842(n1056,n228,n1055);
and gate_843(n1057,n224,n1056);
and gate_844(n1058,n321,n1057);
not gate_845(n1059,n1058);
and gate_846(n1060,n1054,n1059);
and gate_847(n1061,n1045,n1060);
not gate_848(po20,n1061);
and gate_849(n1063,n325,n923);
not gate_850(n1064,n1063);
and gate_851(n1065,pi013,n305);
not gate_852(n1066,n1065);
and gate_853(n1067,pi021,n347);
and gate_854(n1068,n304,n1067);
not gate_855(n1069,n1068);
and gate_856(n1070,n1066,n1069);
and gate_857(n1071,n1064,n1070);
and gate_858(n1072,pi028,n346);
and gate_859(n1073,n304,n1072);
and gate_860(n1074,n324,n1073);
and gate_861(n1075,n333,n1074);
not gate_862(n1076,n1075);
and gate_863(n1077,n351,n1076);
and gate_864(n1078,n1071,n1077);
not gate_865(n1079,n1078);
and gate_866(n1080,n750,n1079);
not gate_867(n1081,n1080);
and gate_868(n1082,n748,n1079);
and gate_869(n1083,n696,n1082);
and gate_870(n1084,pi005,n1083);
not gate_871(n1085,n1084);
and gate_872(n1086,n219,pi115);
and gate_873(n1087,n749,n1086);
and gate_874(n1088,n245,n1087);
not gate_875(n1089,n1088);
and gate_876(n1090,n1085,n1089);
and gate_877(n1091,pi071,n749);
and gate_878(n1092,n228,n1091);
and gate_879(n1093,n224,n1092);
and gate_880(n1094,n321,n1093);
not gate_881(n1095,n1094);
and gate_882(n1096,n1090,n1095);
and gate_883(n1097,n1081,n1096);
not gate_884(po21,n1097);
and gate_885(n1099,n325,n961);
not gate_886(n1100,n1099);
and gate_887(n1101,pi014,n305);
not gate_888(n1102,n1101);
and gate_889(n1103,pi022,n347);
and gate_890(n1104,n304,n1103);
not gate_891(n1105,n1104);
and gate_892(n1106,n1102,n1105);
and gate_893(n1107,n1100,n1106);
and gate_894(n1108,pi029,n346);
and gate_895(n1109,n304,n1108);
and gate_896(n1110,n324,n1109);
and gate_897(n1111,n333,n1110);
not gate_898(n1112,n1111);
and gate_899(n1113,n351,n1112);
and gate_900(n1114,n1107,n1113);
not gate_901(n1115,n1114);
and gate_902(n1116,n750,n1115);
not gate_903(n1117,n1116);
and gate_904(n1118,n748,n1115);
and gate_905(n1119,n696,n1118);
and gate_906(n1120,pi005,n1119);
not gate_907(n1121,n1120);
and gate_908(n1122,n219,pi116);
and gate_909(n1123,n749,n1122);
and gate_910(n1124,n245,n1123);
not gate_911(n1125,n1124);
and gate_912(n1126,n1121,n1125);
and gate_913(n1127,pi072,n749);
and gate_914(n1128,n228,n1127);
and gate_915(n1129,n224,n1128);
and gate_916(n1130,n321,n1129);
not gate_917(n1131,n1130);
and gate_918(n1132,n1126,n1131);
and gate_919(n1133,n1117,n1132);
not gate_920(po22,n1133);
and gate_921(n1135,n325,n999);
not gate_922(n1136,n1135);
and gate_923(n1137,pi015,n305);
not gate_924(n1138,n1137);
and gate_925(n1139,pi023,n347);
and gate_926(n1140,n304,n1139);
not gate_927(n1141,n1140);
and gate_928(n1142,n1138,n1141);
and gate_929(n1143,n1136,n1142);
and gate_930(n1144,pi030,n346);
and gate_931(n1145,n304,n1144);
and gate_932(n1146,n324,n1145);
and gate_933(n1147,n333,n1146);
not gate_934(n1148,n1147);
and gate_935(n1149,n351,n1148);
and gate_936(n1150,n1143,n1149);
not gate_937(n1151,n1150);
and gate_938(n1152,n750,n1151);
not gate_939(n1153,n1152);
and gate_940(n1154,n748,n1151);
and gate_941(n1155,n696,n1154);
and gate_942(n1156,pi005,n1155);
not gate_943(n1157,n1156);
and gate_944(n1158,n219,pi117);
and gate_945(n1159,n749,n1158);
and gate_946(n1160,n245,n1159);
not gate_947(n1161,n1160);
and gate_948(n1162,n1157,n1161);
and gate_949(n1163,pi073,n749);
and gate_950(n1164,n228,n1163);
and gate_951(n1165,n224,n1164);
and gate_952(n1166,n321,n1165);
not gate_953(n1167,n1166);
and gate_954(n1168,n1162,n1167);
and gate_955(n1169,n1153,n1168);
not gate_956(po23,n1169);
and gate_957(n1171,n325,n1037);
not gate_958(n1172,n1171);
and gate_959(n1173,pi016,n305);
not gate_960(n1174,n1173);
and gate_961(n1175,pi024,n347);
and gate_962(n1176,n304,n1175);
not gate_963(n1177,n1176);
and gate_964(n1178,n1174,n1177);
and gate_965(n1179,n1172,n1178);
and gate_966(n1180,pi031,n346);
and gate_967(n1181,n304,n1180);
and gate_968(n1182,n324,n1181);
and gate_969(n1183,n333,n1182);
not gate_970(n1184,n1183);
and gate_971(n1185,n351,n1184);
and gate_972(n1186,n1179,n1185);
not gate_973(n1187,n1186);
and gate_974(n1188,n750,n1187);
not gate_975(n1189,n1188);
and gate_976(n1190,n748,n1187);
and gate_977(n1191,n696,n1190);
and gate_978(n1192,pi005,n1191);
not gate_979(n1193,n1192);
and gate_980(n1194,n219,pi118);
and gate_981(n1195,n749,n1194);
and gate_982(n1196,n245,n1195);
not gate_983(n1197,n1196);
and gate_984(n1198,n1193,n1197);
and gate_985(n1199,pi074,n749);
and gate_986(n1200,n228,n1199);
and gate_987(n1201,n224,n1200);
and gate_988(n1202,n321,n1201);
not gate_989(n1203,n1202);
and gate_990(n1204,n1198,n1203);
and gate_991(n1205,n1189,n1204);
not gate_992(po24,n1205);
and gate_993(n1207,n325,n1073);
not gate_994(n1208,n1207);
and gate_995(n1209,pi017,n305);
not gate_996(n1210,n1209);
and gate_997(n1211,pi025,n347);
and gate_998(n1212,n304,n1211);
not gate_999(n1213,n1212);
and gate_1000(n1214,n1210,n1213);
and gate_1001(n1215,n1208,n1214);
and gate_1002(n1216,pi032,n346);
and gate_1003(n1217,n304,n1216);
and gate_1004(n1218,n324,n1217);
and gate_1005(n1219,n333,n1218);
not gate_1006(n1220,n1219);
and gate_1007(n1221,n351,n1220);
and gate_1008(n1222,n1215,n1221);
not gate_1009(n1223,n1222);
and gate_1010(n1224,n750,n1223);
not gate_1011(n1225,n1224);
and gate_1012(n1226,n748,n1223);
and gate_1013(n1227,n696,n1226);
and gate_1014(n1228,pi005,n1227);
not gate_1015(n1229,n1228);
and gate_1016(n1230,n219,pi119);
and gate_1017(n1231,n749,n1230);
and gate_1018(n1232,n245,n1231);
not gate_1019(n1233,n1232);
and gate_1020(n1234,n1229,n1233);
and gate_1021(n1235,pi075,n749);
and gate_1022(n1236,n228,n1235);
and gate_1023(n1237,n224,n1236);
and gate_1024(n1238,n321,n1237);
not gate_1025(n1239,n1238);
and gate_1026(n1240,n1234,n1239);
and gate_1027(n1241,n1225,n1240);
not gate_1028(po25,n1241);
and gate_1029(n1243,n325,n1109);
not gate_1030(n1244,n1243);
and gate_1031(n1245,pi018,n305);
not gate_1032(n1246,n1245);
and gate_1033(n1247,pi026,n347);
and gate_1034(n1248,n304,n1247);
not gate_1035(n1249,n1248);
and gate_1036(n1250,n1246,n1249);
and gate_1037(n1251,n1244,n1250);
and gate_1038(n1252,pi033,n346);
and gate_1039(n1253,n304,n1252);
and gate_1040(n1254,n324,n1253);
and gate_1041(n1255,n333,n1254);
not gate_1042(n1256,n1255);
and gate_1043(n1257,n351,n1256);
and gate_1044(n1258,n1251,n1257);
not gate_1045(n1259,n1258);
and gate_1046(n1260,n750,n1259);
not gate_1047(n1261,n1260);
and gate_1048(n1262,n748,n1259);
and gate_1049(n1263,n696,n1262);
and gate_1050(n1264,pi005,n1263);
not gate_1051(n1265,n1264);
and gate_1052(n1266,n219,pi120);
and gate_1053(n1267,n749,n1266);
and gate_1054(n1268,n245,n1267);
not gate_1055(n1269,n1268);
and gate_1056(n1270,n1265,n1269);
and gate_1057(n1271,pi076,n749);
and gate_1058(n1272,n228,n1271);
and gate_1059(n1273,n224,n1272);
and gate_1060(n1274,n321,n1273);
not gate_1061(n1275,n1274);
and gate_1062(n1276,n1270,n1275);
and gate_1063(n1277,n1261,n1276);
not gate_1064(po26,n1277);
and gate_1065(n1279,n325,n1145);
not gate_1066(n1280,n1279);
and gate_1067(n1281,pi019,n305);
not gate_1068(n1282,n1281);
and gate_1069(n1283,pi027,n347);
and gate_1070(n1284,n304,n1283);
not gate_1071(n1285,n1284);
and gate_1072(n1286,n1282,n1285);
and gate_1073(n1287,n1280,n1286);
and gate_1074(n1288,pi034,n346);
and gate_1075(n1289,n304,n1288);
and gate_1076(n1290,n324,n1289);
and gate_1077(n1291,n333,n1290);
not gate_1078(n1292,n1291);
and gate_1079(n1293,n351,n1292);
and gate_1080(n1294,n1287,n1293);
not gate_1081(n1295,n1294);
and gate_1082(n1296,n750,n1295);
not gate_1083(n1297,n1296);
and gate_1084(n1298,n748,n1295);
and gate_1085(n1299,n696,n1298);
and gate_1086(n1300,pi005,n1299);
not gate_1087(n1301,n1300);
and gate_1088(n1302,n219,pi121);
and gate_1089(n1303,n749,n1302);
and gate_1090(n1304,n245,n1303);
not gate_1091(n1305,n1304);
and gate_1092(n1306,n1301,n1305);
and gate_1093(n1307,pi077,n749);
and gate_1094(n1308,n228,n1307);
and gate_1095(n1309,n224,n1308);
and gate_1096(n1310,n321,n1309);
not gate_1097(n1311,n1310);
and gate_1098(n1312,n1306,n1311);
and gate_1099(n1313,n1297,n1312);
not gate_1100(po27,n1313);
and gate_1101(n1315,n325,n1181);
not gate_1102(n1316,n1315);
and gate_1103(n1317,pi020,n305);
not gate_1104(n1318,n1317);
and gate_1105(n1319,pi028,n347);
and gate_1106(n1320,n304,n1319);
not gate_1107(n1321,n1320);
and gate_1108(n1322,n1318,n1321);
and gate_1109(n1323,n1316,n1322);
and gate_1110(n1324,n324,n857);
and gate_1111(n1325,n333,n1324);
not gate_1112(n1326,n1325);
and gate_1113(n1327,n351,n1326);
and gate_1114(n1328,n1323,n1327);
not gate_1115(n1329,n1328);
and gate_1116(n1330,n750,n1329);
not gate_1117(n1331,n1330);
and gate_1118(n1332,n748,n1329);
and gate_1119(n1333,n696,n1332);
and gate_1120(n1334,pi005,n1333);
not gate_1121(n1335,n1334);
and gate_1122(n1336,n219,pi122);
and gate_1123(n1337,n749,n1336);
and gate_1124(n1338,n245,n1337);
not gate_1125(n1339,n1338);
and gate_1126(n1340,n1335,n1339);
and gate_1127(n1341,pi078,n749);
and gate_1128(n1342,n228,n1341);
and gate_1129(n1343,n224,n1342);
and gate_1130(n1344,n321,n1343);
not gate_1131(n1345,n1344);
and gate_1132(n1346,n1340,n1345);
and gate_1133(n1347,n1331,n1346);
not gate_1134(po28,n1347);
and gate_1135(n1349,n325,n1217);
not gate_1136(n1350,n1349);
and gate_1137(n1351,pi021,n305);
not gate_1138(n1352,n1351);
and gate_1139(n1353,pi029,n347);
and gate_1140(n1354,n304,n1353);
not gate_1141(n1355,n1354);
and gate_1142(n1356,n1352,n1355);
and gate_1143(n1357,n1350,n1356);
and gate_1144(n1358,n324,n727);
and gate_1145(n1359,n333,n1358);
not gate_1146(n1360,n1359);
and gate_1147(n1361,n351,n1360);
and gate_1148(n1362,n1357,n1361);
not gate_1149(n1363,n1362);
and gate_1150(n1364,n750,n1363);
not gate_1151(n1365,n1364);
and gate_1152(n1366,n748,n1363);
and gate_1153(n1367,n696,n1366);
and gate_1154(n1368,pi005,n1367);
not gate_1155(n1369,n1368);
and gate_1156(n1370,n219,pi123);
and gate_1157(n1371,n749,n1370);
and gate_1158(n1372,n245,n1371);
not gate_1159(n1373,n1372);
and gate_1160(n1374,n1369,n1373);
and gate_1161(n1375,pi079,n749);
and gate_1162(n1376,n228,n1375);
and gate_1163(n1377,n224,n1376);
and gate_1164(n1378,n321,n1377);
not gate_1165(n1379,n1378);
and gate_1166(n1380,n1374,n1379);
and gate_1167(n1381,n1365,n1380);
not gate_1168(po29,n1381);
and gate_1169(n1383,n325,n1253);
not gate_1170(n1384,n1383);
and gate_1171(n1385,pi022,n305);
not gate_1172(n1386,n1385);
and gate_1173(n1387,pi030,n347);
and gate_1174(n1388,n304,n1387);
not gate_1175(n1389,n1388);
and gate_1176(n1390,n1386,n1389);
and gate_1177(n1391,n1384,n1390);
and gate_1178(n1392,n324,n778);
and gate_1179(n1393,n333,n1392);
not gate_1180(n1394,n1393);
and gate_1181(n1395,n351,n1394);
and gate_1182(n1396,n1391,n1395);
not gate_1183(n1397,n1396);
and gate_1184(n1398,n750,n1397);
not gate_1185(n1399,n1398);
and gate_1186(n1400,n748,n1397);
and gate_1187(n1401,n696,n1400);
and gate_1188(n1402,pi005,n1401);
not gate_1189(n1403,n1402);
and gate_1190(n1404,n219,pi124);
and gate_1191(n1405,n749,n1404);
and gate_1192(n1406,n245,n1405);
not gate_1193(n1407,n1406);
and gate_1194(n1408,n1403,n1407);
and gate_1195(n1409,pi080,n749);
and gate_1196(n1410,n228,n1409);
and gate_1197(n1411,n224,n1410);
and gate_1198(n1412,n321,n1411);
not gate_1199(n1413,n1412);
and gate_1200(n1414,n1408,n1413);
and gate_1201(n1415,n1399,n1414);
not gate_1202(po30,n1415);
and gate_1203(n1417,n325,n1289);
not gate_1204(n1418,n1417);
and gate_1205(n1419,pi023,n305);
not gate_1206(n1420,n1419);
and gate_1207(n1421,pi031,n347);
and gate_1208(n1422,n304,n1421);
not gate_1209(n1423,n1422);
and gate_1210(n1424,n1420,n1423);
and gate_1211(n1425,n1418,n1424);
and gate_1212(n1426,n324,n816);
and gate_1213(n1427,n333,n1426);
not gate_1214(n1428,n1427);
and gate_1215(n1429,n351,n1428);
and gate_1216(n1430,n1425,n1429);
not gate_1217(n1431,n1430);
and gate_1218(n1432,n750,n1431);
not gate_1219(n1433,n1432);
and gate_1220(n1434,n748,n1431);
and gate_1221(n1435,n696,n1434);
and gate_1222(n1436,pi005,n1435);
not gate_1223(n1437,n1436);
and gate_1224(n1438,n219,pi125);
and gate_1225(n1439,n749,n1438);
and gate_1226(n1440,n245,n1439);
not gate_1227(n1441,n1440);
and gate_1228(n1442,n1437,n1441);
and gate_1229(n1443,pi081,n749);
and gate_1230(n1444,n228,n1443);
and gate_1231(n1445,n224,n1444);
and gate_1232(n1446,n321,n1445);
not gate_1233(n1447,n1446);
and gate_1234(n1448,n1442,n1447);
and gate_1235(n1449,n1433,n1448);
not gate_1236(po31,n1449);
and gate_1237(n1451,pi007,n688);
not gate_1238(n1452,n1451);
and gate_1239(n1453,pi000,n274);
and gate_1240(n1454,n224,n1453);
and gate_1241(n1455,n220,n1454);
not gate_1242(n1456,n1455);
and gate_1243(n1457,pi078,n346);
and gate_1244(n1458,n304,n1457);
and gate_1245(n1459,n325,n1458);
not gate_1246(n1460,n1459);
and gate_1247(n1461,pi067,n305);
not gate_1248(n1462,n1461);
and gate_1249(n1463,pi075,n347);
and gate_1250(n1464,n304,n1463);
not gate_1251(n1465,n1464);
and gate_1252(n1466,n1462,n1465);
and gate_1253(n1467,n1460,n1466);
and gate_1254(n1468,pi082,n346);
and gate_1255(n1469,n304,n1468);
and gate_1256(n1470,n324,n1469);
and gate_1257(n1471,n333,n1470);
not gate_1258(n1472,n1471);
and gate_1259(n1473,n351,n1472);
and gate_1260(n1474,n1467,n1473);
not gate_1261(n1475,n1474);
and gate_1262(n1476,pi003,n225);
and gate_1263(n1477,n688,n1476);
and gate_1264(n1478,pi004,n1477);
not gate_1265(n1479,n1478);
and gate_1266(n1480,n1475,n1479);
and gate_1267(n1481,n218,n746);
not gate_1268(n1482,n1481);
and gate_1269(n1483,n1480,n1482);
and gate_1270(n1484,n217,pi004);
and gate_1271(n1485,n688,n1484);
not gate_1272(n1486,n1485);
and gate_1273(n1487,n1483,n1486);
and gate_1274(n1488,n1456,n1487);
and gate_1275(n1489,n1451,n1488);
not gate_1276(n1490,n1489);
and gate_1277(n1491,n1452,n1475);
and gate_1278(n1492,n1486,n1491);
and gate_1279(n1493,n1482,n1492);
and gate_1280(n1494,n1479,n1493);
and gate_1281(n1495,n1456,n1494);
and gate_1282(n1496,pi005,n1495);
not gate_1283(n1497,n1496);
and gate_1284(n1498,n1490,n1497);
and gate_1285(n1499,n936,n1456);
and gate_1286(n1500,n1479,n1499);
and gate_1287(n1501,n1482,n1500);
and gate_1288(n1502,n1486,n1501);
and gate_1289(n1503,n245,n1502);
not gate_1290(n1504,n1503);
and gate_1291(n1505,n1498,n1504);
and gate_1292(n1506,n1479,n1482);
and gate_1293(n1507,n1456,n1486);
and gate_1294(n1508,n1506,n1507);
not gate_1295(n1509,n1508);
and gate_1296(n1510,n1475,n1509);
not gate_1297(n1511,n1510);
and gate_1298(n1512,n1505,n1511);
not gate_1299(po32,n1512);
and gate_1300(n1514,pi079,n346);
and gate_1301(n1515,n304,n1514);
and gate_1302(n1516,n325,n1515);
not gate_1303(n1517,n1516);
and gate_1304(n1518,pi068,n305);
not gate_1305(n1519,n1518);
and gate_1306(n1520,pi076,n347);
and gate_1307(n1521,n304,n1520);
not gate_1308(n1522,n1521);
and gate_1309(n1523,n1519,n1522);
and gate_1310(n1524,n1517,n1523);
and gate_1311(n1525,pi083,n346);
and gate_1312(n1526,n304,n1525);
and gate_1313(n1527,n324,n1526);
and gate_1314(n1528,n333,n1527);
not gate_1315(n1529,n1528);
and gate_1316(n1530,n351,n1529);
and gate_1317(n1531,n1524,n1530);
not gate_1318(n1532,n1531);
and gate_1319(n1533,n1506,n1532);
and gate_1320(n1534,n1507,n1533);
and gate_1321(n1535,n1451,n1534);
not gate_1322(n1536,n1535);
and gate_1323(n1537,n1452,n1532);
and gate_1324(n1538,n1508,n1537);
and gate_1325(n1539,pi005,n1538);
not gate_1326(n1540,n1539);
and gate_1327(n1541,n1536,n1540);
and gate_1328(n1542,n974,n1508);
and gate_1329(n1543,n245,n1542);
not gate_1330(n1544,n1543);
and gate_1331(n1545,n1541,n1544);
and gate_1332(n1546,n1509,n1532);
not gate_1333(n1547,n1546);
and gate_1334(n1548,n1545,n1547);
not gate_1335(po33,n1548);
and gate_1336(n1550,pi080,n346);
and gate_1337(n1551,n304,n1550);
and gate_1338(n1552,n325,n1551);
not gate_1339(n1553,n1552);
and gate_1340(n1554,pi069,n305);
not gate_1341(n1555,n1554);
and gate_1342(n1556,pi077,n347);
and gate_1343(n1557,n304,n1556);
not gate_1344(n1558,n1557);
and gate_1345(n1559,n1555,n1558);
and gate_1346(n1560,n1553,n1559);
and gate_1347(n1561,pi084,n346);
and gate_1348(n1562,n304,n1561);
and gate_1349(n1563,n324,n1562);
and gate_1350(n1564,n333,n1563);
not gate_1351(n1565,n1564);
and gate_1352(n1566,n351,n1565);
and gate_1353(n1567,n1560,n1566);
not gate_1354(n1568,n1567);
and gate_1355(n1569,n1506,n1568);
and gate_1356(n1570,n1507,n1569);
and gate_1357(n1571,n1451,n1570);
not gate_1358(n1572,n1571);
and gate_1359(n1573,n1452,n1568);
and gate_1360(n1574,n1508,n1573);
and gate_1361(n1575,pi005,n1574);
not gate_1362(n1576,n1575);
and gate_1363(n1577,n1572,n1576);
and gate_1364(n1578,n1012,n1508);
and gate_1365(n1579,n245,n1578);
not gate_1366(n1580,n1579);
and gate_1367(n1581,n1577,n1580);
and gate_1368(n1582,n1509,n1568);
not gate_1369(n1583,n1582);
and gate_1370(n1584,n1581,n1583);
not gate_1371(po34,n1584);
and gate_1372(n1586,pi081,n346);
and gate_1373(n1587,n304,n1586);
and gate_1374(n1588,n325,n1587);
not gate_1375(n1589,n1588);
and gate_1376(n1590,pi070,n305);
not gate_1377(n1591,n1590);
and gate_1378(n1592,pi078,n347);
and gate_1379(n1593,n304,n1592);
not gate_1380(n1594,n1593);
and gate_1381(n1595,n1591,n1594);
and gate_1382(n1596,n1589,n1595);
and gate_1383(n1597,pi085,n346);
and gate_1384(n1598,n304,n1597);
and gate_1385(n1599,n324,n1598);
and gate_1386(n1600,n333,n1599);
not gate_1387(n1601,n1600);
and gate_1388(n1602,n351,n1601);
and gate_1389(n1603,n1596,n1602);
not gate_1390(n1604,n1603);
and gate_1391(n1605,n1506,n1604);
and gate_1392(n1606,n1507,n1605);
and gate_1393(n1607,n1451,n1606);
not gate_1394(n1608,n1607);
and gate_1395(n1609,n1452,n1604);
and gate_1396(n1610,n1508,n1609);
and gate_1397(n1611,pi005,n1610);
not gate_1398(n1612,n1611);
and gate_1399(n1613,n1608,n1612);
and gate_1400(n1614,n1050,n1508);
and gate_1401(n1615,n245,n1614);
not gate_1402(n1616,n1615);
and gate_1403(n1617,n1613,n1616);
and gate_1404(n1618,n1509,n1604);
not gate_1405(n1619,n1618);
and gate_1406(n1620,n1617,n1619);
not gate_1407(po35,n1620);
and gate_1408(n1622,n325,n1469);
not gate_1409(n1623,n1622);
and gate_1410(n1624,pi071,n305);
not gate_1411(n1625,n1624);
and gate_1412(n1626,pi079,n347);
and gate_1413(n1627,n304,n1626);
not gate_1414(n1628,n1627);
and gate_1415(n1629,n1625,n1628);
and gate_1416(n1630,n1623,n1629);
and gate_1417(n1631,pi086,n346);
and gate_1418(n1632,n304,n1631);
and gate_1419(n1633,n324,n1632);
and gate_1420(n1634,n333,n1633);
not gate_1421(n1635,n1634);
and gate_1422(n1636,n351,n1635);
and gate_1423(n1637,n1630,n1636);
not gate_1424(n1638,n1637);
and gate_1425(n1639,n1506,n1638);
and gate_1426(n1640,n1507,n1639);
and gate_1427(n1641,n1451,n1640);
not gate_1428(n1642,n1641);
and gate_1429(n1643,n1452,n1638);
and gate_1430(n1644,n1508,n1643);
and gate_1431(n1645,pi005,n1644);
not gate_1432(n1646,n1645);
and gate_1433(n1647,n1642,n1646);
and gate_1434(n1648,n1086,n1508);
and gate_1435(n1649,n245,n1648);
not gate_1436(n1650,n1649);
and gate_1437(n1651,n1647,n1650);
and gate_1438(n1652,n1509,n1638);
not gate_1439(n1653,n1652);
and gate_1440(n1654,n1651,n1653);
not gate_1441(po36,n1654);
and gate_1442(n1656,n325,n1526);
not gate_1443(n1657,n1656);
and gate_1444(n1658,pi072,n305);
not gate_1445(n1659,n1658);
and gate_1446(n1660,pi080,n347);
and gate_1447(n1661,n304,n1660);
not gate_1448(n1662,n1661);
and gate_1449(n1663,n1659,n1662);
and gate_1450(n1664,n1657,n1663);
and gate_1451(n1665,n324,n619);
and gate_1452(n1666,n333,n1665);
not gate_1453(n1667,n1666);
and gate_1454(n1668,n351,n1667);
and gate_1455(n1669,n1664,n1668);
not gate_1456(n1670,n1669);
and gate_1457(n1671,n1506,n1670);
and gate_1458(n1672,n1507,n1671);
and gate_1459(n1673,n1451,n1672);
not gate_1460(n1674,n1673);
and gate_1461(n1675,n1452,n1670);
and gate_1462(n1676,n1508,n1675);
and gate_1463(n1677,pi005,n1676);
not gate_1464(n1678,n1677);
and gate_1465(n1679,n1674,n1678);
and gate_1466(n1680,n1122,n1508);
and gate_1467(n1681,n245,n1680);
not gate_1468(n1682,n1681);
and gate_1469(n1683,n1679,n1682);
and gate_1470(n1684,n1509,n1670);
not gate_1471(n1685,n1684);
and gate_1472(n1686,n1683,n1685);
not gate_1473(po37,n1686);
and gate_1474(n1688,n325,n1562);
not gate_1475(n1689,n1688);
and gate_1476(n1690,pi073,n305);
not gate_1477(n1691,n1690);
and gate_1478(n1692,pi081,n347);
and gate_1479(n1693,n304,n1692);
not gate_1480(n1694,n1693);
and gate_1481(n1695,n1691,n1694);
and gate_1482(n1696,n1689,n1695);
and gate_1483(n1697,n324,n647);
and gate_1484(n1698,n333,n1697);
not gate_1485(n1699,n1698);
and gate_1486(n1700,n351,n1699);
and gate_1487(n1701,n1696,n1700);
not gate_1488(n1702,n1701);
and gate_1489(n1703,n1506,n1702);
and gate_1490(n1704,n1507,n1703);
and gate_1491(n1705,n1451,n1704);
not gate_1492(n1706,n1705);
and gate_1493(n1707,n1452,n1702);
and gate_1494(n1708,n1508,n1707);
and gate_1495(n1709,pi005,n1708);
not gate_1496(n1710,n1709);
and gate_1497(n1711,n1706,n1710);
and gate_1498(n1712,n1158,n1508);
and gate_1499(n1713,n245,n1712);
not gate_1500(n1714,n1713);
and gate_1501(n1715,n1711,n1714);
and gate_1502(n1716,n1509,n1702);
not gate_1503(n1717,n1716);
and gate_1504(n1718,n1715,n1717);
not gate_1505(po38,n1718);
and gate_1506(n1720,n325,n1598);
not gate_1507(n1721,n1720);
and gate_1508(n1722,pi074,n305);
not gate_1509(n1723,n1722);
and gate_1510(n1724,pi082,n347);
and gate_1511(n1725,n304,n1724);
not gate_1512(n1726,n1725);
and gate_1513(n1727,n1723,n1726);
and gate_1514(n1728,n1721,n1727);
and gate_1515(n1729,n324,n580);
and gate_1516(n1730,n333,n1729);
not gate_1517(n1731,n1730);
and gate_1518(n1732,n351,n1731);
and gate_1519(n1733,n1728,n1732);
not gate_1520(n1734,n1733);
and gate_1521(n1735,n1506,n1734);
and gate_1522(n1736,n1507,n1735);
and gate_1523(n1737,n1451,n1736);
not gate_1524(n1738,n1737);
and gate_1525(n1739,n1452,n1734);
and gate_1526(n1740,n1508,n1739);
and gate_1527(n1741,pi005,n1740);
not gate_1528(n1742,n1741);
and gate_1529(n1743,n1738,n1742);
and gate_1530(n1744,n1194,n1508);
and gate_1531(n1745,n245,n1744);
not gate_1532(n1746,n1745);
and gate_1533(n1747,n1743,n1746);
and gate_1534(n1748,n1509,n1734);
not gate_1535(n1749,n1748);
and gate_1536(n1750,n1747,n1749);
not gate_1537(po39,n1750);
and gate_1538(n1752,n325,n1632);
not gate_1539(n1753,n1752);
and gate_1540(n1754,pi075,n305);
not gate_1541(n1755,n1754);
and gate_1542(n1756,pi083,n347);
and gate_1543(n1757,n304,n1756);
not gate_1544(n1758,n1757);
and gate_1545(n1759,n1755,n1758);
and gate_1546(n1760,n1753,n1759);
and gate_1547(n1761,n324,n423);
and gate_1548(n1762,n333,n1761);
not gate_1549(n1763,n1762);
and gate_1550(n1764,n351,n1763);
and gate_1551(n1765,n1760,n1764);
not gate_1552(n1766,n1765);
and gate_1553(n1767,n1506,n1766);
and gate_1554(n1768,n1507,n1767);
and gate_1555(n1769,n1451,n1768);
not gate_1556(n1770,n1769);
and gate_1557(n1771,n1452,n1766);
and gate_1558(n1772,n1508,n1771);
and gate_1559(n1773,pi005,n1772);
not gate_1560(n1774,n1773);
and gate_1561(n1775,n1770,n1774);
and gate_1562(n1776,n1230,n1508);
and gate_1563(n1777,n245,n1776);
not gate_1564(n1778,n1777);
and gate_1565(n1779,n1775,n1778);
and gate_1566(n1780,n1509,n1766);
not gate_1567(n1781,n1780);
and gate_1568(n1782,n1779,n1781);
not gate_1569(po40,n1782);
and gate_1570(n1784,pi076,n305);
not gate_1571(n1785,n1784);
and gate_1572(n1786,pi084,n347);
and gate_1573(n1787,n304,n1786);
not gate_1574(n1788,n1787);
and gate_1575(n1789,n1785,n1788);
and gate_1576(n1790,n621,n1789);
and gate_1577(n1791,n324,n466);
and gate_1578(n1792,n333,n1791);
not gate_1579(n1793,n1792);
and gate_1580(n1794,n351,n1793);
and gate_1581(n1795,n1790,n1794);
not gate_1582(n1796,n1795);
and gate_1583(n1797,n1506,n1796);
and gate_1584(n1798,n1507,n1797);
and gate_1585(n1799,n1451,n1798);
not gate_1586(n1800,n1799);
and gate_1587(n1801,n1452,n1796);
and gate_1588(n1802,n1508,n1801);
and gate_1589(n1803,pi005,n1802);
not gate_1590(n1804,n1803);
and gate_1591(n1805,n1800,n1804);
and gate_1592(n1806,n1266,n1508);
and gate_1593(n1807,n245,n1806);
not gate_1594(n1808,n1807);
and gate_1595(n1809,n1805,n1808);
and gate_1596(n1810,n1509,n1796);
not gate_1597(n1811,n1810);
and gate_1598(n1812,n1809,n1811);
not gate_1599(po41,n1812);
and gate_1600(n1814,pi077,n305);
not gate_1601(n1815,n1814);
and gate_1602(n1816,pi085,n347);
and gate_1603(n1817,n304,n1816);
not gate_1604(n1818,n1817);
and gate_1605(n1819,n1815,n1818);
and gate_1606(n1820,n649,n1819);
and gate_1607(n1821,n324,n492);
and gate_1608(n1822,n333,n1821);
not gate_1609(n1823,n1822);
and gate_1610(n1824,n351,n1823);
and gate_1611(n1825,n1820,n1824);
not gate_1612(n1826,n1825);
and gate_1613(n1827,n1506,n1826);
and gate_1614(n1828,n1507,n1827);
and gate_1615(n1829,n1451,n1828);
not gate_1616(n1830,n1829);
and gate_1617(n1831,n1452,n1826);
and gate_1618(n1832,n1508,n1831);
and gate_1619(n1833,pi005,n1832);
not gate_1620(n1834,n1833);
and gate_1621(n1835,n1830,n1834);
and gate_1622(n1836,n1302,n1508);
and gate_1623(n1837,n245,n1836);
not gate_1624(n1838,n1837);
and gate_1625(n1839,n1835,n1838);
and gate_1626(n1840,n1509,n1826);
not gate_1627(n1841,n1840);
and gate_1628(n1842,n1839,n1841);
not gate_1629(po42,n1842);
and gate_1630(n1844,pi078,n305);
not gate_1631(n1845,n1844);
and gate_1632(n1846,pi086,n347);
and gate_1633(n1847,n304,n1846);
not gate_1634(n1848,n1847);
and gate_1635(n1849,n1845,n1848);
and gate_1636(n1850,n582,n1849);
and gate_1637(n1851,n324,n516);
and gate_1638(n1852,n333,n1851);
not gate_1639(n1853,n1852);
and gate_1640(n1854,n351,n1853);
and gate_1641(n1855,n1850,n1854);
not gate_1642(n1856,n1855);
and gate_1643(n1857,n1506,n1856);
and gate_1644(n1858,n1507,n1857);
and gate_1645(n1859,n1451,n1858);
not gate_1646(n1860,n1859);
and gate_1647(n1861,n1452,n1856);
and gate_1648(n1862,n1508,n1861);
and gate_1649(n1863,pi005,n1862);
not gate_1650(n1864,n1863);
and gate_1651(n1865,n1860,n1864);
and gate_1652(n1866,n1336,n1508);
and gate_1653(n1867,n245,n1866);
not gate_1654(n1868,n1867);
and gate_1655(n1869,n1865,n1868);
and gate_1656(n1870,n1509,n1856);
not gate_1657(n1871,n1870);
and gate_1658(n1872,n1869,n1871);
not gate_1659(po43,n1872);
and gate_1660(n1874,pi079,n305);
not gate_1661(n1875,n1874);
and gate_1662(n1876,pi041,n347);
and gate_1663(n1877,n304,n1876);
not gate_1664(n1878,n1877);
and gate_1665(n1879,n1875,n1878);
and gate_1666(n1880,n425,n1879);
and gate_1667(n1881,n324,n540);
and gate_1668(n1882,n333,n1881);
not gate_1669(n1883,n1882);
and gate_1670(n1884,n351,n1883);
and gate_1671(n1885,n1880,n1884);
not gate_1672(n1886,n1885);
and gate_1673(n1887,n1506,n1886);
and gate_1674(n1888,n1507,n1887);
and gate_1675(n1889,n1451,n1888);
not gate_1676(n1890,n1889);
and gate_1677(n1891,n1452,n1886);
and gate_1678(n1892,n1508,n1891);
and gate_1679(n1893,pi005,n1892);
not gate_1680(n1894,n1893);
and gate_1681(n1895,n1890,n1894);
and gate_1682(n1896,n1370,n1508);
and gate_1683(n1897,n245,n1896);
not gate_1684(n1898,n1897);
and gate_1685(n1899,n1895,n1898);
and gate_1686(n1900,n1509,n1886);
not gate_1687(n1901,n1900);
and gate_1688(n1902,n1899,n1901);
not gate_1689(po44,n1902);
and gate_1690(n1904,pi080,n305);
not gate_1691(n1905,n1904);
and gate_1692(n1906,pi042,n347);
and gate_1693(n1907,n304,n1906);
not gate_1694(n1908,n1907);
and gate_1695(n1909,n1905,n1908);
and gate_1696(n1910,n468,n1909);
and gate_1697(n1911,n324,n564);
and gate_1698(n1912,n333,n1911);
not gate_1699(n1913,n1912);
and gate_1700(n1914,n351,n1913);
and gate_1701(n1915,n1910,n1914);
not gate_1702(n1916,n1915);
and gate_1703(n1917,n1506,n1916);
and gate_1704(n1918,n1507,n1917);
and gate_1705(n1919,n1451,n1918);
not gate_1706(n1920,n1919);
and gate_1707(n1921,n1452,n1916);
and gate_1708(n1922,n1508,n1921);
and gate_1709(n1923,pi005,n1922);
not gate_1710(n1924,n1923);
and gate_1711(n1925,n1920,n1924);
and gate_1712(n1926,n1404,n1508);
and gate_1713(n1927,n245,n1926);
not gate_1714(n1928,n1927);
and gate_1715(n1929,n1925,n1928);
and gate_1716(n1930,n1509,n1916);
not gate_1717(n1931,n1930);
and gate_1718(n1932,n1929,n1931);
not gate_1719(po45,n1932);
and gate_1720(n1934,pi081,n305);
not gate_1721(n1935,n1934);
and gate_1722(n1936,pi043,n347);
and gate_1723(n1937,n304,n1936);
not gate_1724(n1938,n1937);
and gate_1725(n1939,n1935,n1938);
and gate_1726(n1940,n494,n1939);
and gate_1727(n1941,n324,n354);
and gate_1728(n1942,n333,n1941);
not gate_1729(n1943,n1942);
and gate_1730(n1944,n351,n1943);
and gate_1731(n1945,n1940,n1944);
not gate_1732(n1946,n1945);
and gate_1733(n1947,n1506,n1946);
and gate_1734(n1948,n1507,n1947);
and gate_1735(n1949,n1451,n1948);
not gate_1736(n1950,n1949);
and gate_1737(n1951,n1452,n1946);
and gate_1738(n1952,n1508,n1951);
and gate_1739(n1953,pi005,n1952);
not gate_1740(n1954,n1953);
and gate_1741(n1955,n1950,n1954);
and gate_1742(n1956,n1438,n1508);
and gate_1743(n1957,n245,n1956);
not gate_1744(n1958,n1957);
and gate_1745(n1959,n1955,n1958);
and gate_1746(n1960,n1509,n1946);
not gate_1747(n1961,n1960);
and gate_1748(n1962,n1959,n1961);
not gate_1749(po46,n1962);
and gate_1750(n1964,pi082,n305);
not gate_1751(n1965,n1964);
and gate_1752(n1966,pi044,n347);
and gate_1753(n1967,n304,n1966);
not gate_1754(n1968,n1967);
and gate_1755(n1969,n1965,n1968);
and gate_1756(n1970,n518,n1969);
and gate_1757(n1971,n324,n376);
and gate_1758(n1972,n333,n1971);
not gate_1759(n1973,n1972);
and gate_1760(n1974,n351,n1973);
and gate_1761(n1975,n1970,n1974);
not gate_1762(n1976,n1975);
and gate_1763(n1977,n1506,n1976);
and gate_1764(n1978,n1507,n1977);
and gate_1765(n1979,n1451,n1978);
not gate_1766(n1980,n1979);
and gate_1767(n1981,n1452,n1976);
and gate_1768(n1982,n1508,n1981);
and gate_1769(n1983,pi005,n1982);
not gate_1770(n1984,n1983);
and gate_1771(n1985,n1980,n1984);
and gate_1772(n1986,n886,n1508);
and gate_1773(n1987,n245,n1986);
not gate_1774(n1988,n1987);
and gate_1775(n1989,n1985,n1988);
and gate_1776(n1990,n1509,n1976);
not gate_1777(n1991,n1990);
and gate_1778(n1992,n1989,n1991);
not gate_1779(po47,n1992);
and gate_1780(n1994,pi083,n305);
not gate_1781(n1995,n1994);
and gate_1782(n1996,pi045,n347);
and gate_1783(n1997,n304,n1996);
not gate_1784(n1998,n1997);
and gate_1785(n1999,n1995,n1998);
and gate_1786(n2000,n542,n1999);
and gate_1787(n2001,pi087,n346);
and gate_1788(n2002,n304,n2001);
and gate_1789(n2003,n324,n2002);
and gate_1790(n2004,n333,n2003);
not gate_1791(n2005,n2004);
and gate_1792(n2006,n351,n2005);
and gate_1793(n2007,n2000,n2006);
not gate_1794(n2008,n2007);
and gate_1795(n2009,n1506,n2008);
and gate_1796(n2010,n1507,n2009);
and gate_1797(n2011,n1451,n2010);
not gate_1798(n2012,n2011);
and gate_1799(n2013,n1452,n2008);
and gate_1800(n2014,n1508,n2013);
and gate_1801(n2015,pi005,n2014);
not gate_1802(n2016,n2015);
and gate_1803(n2017,n2012,n2016);
and gate_1804(n2018,n758,n1508);
and gate_1805(n2019,n245,n2018);
not gate_1806(n2020,n2019);
and gate_1807(n2021,n2017,n2020);
and gate_1808(n2022,n1509,n2008);
not gate_1809(n2023,n2022);
and gate_1810(n2024,n2021,n2023);
not gate_1811(po48,n2024);
and gate_1812(n2026,pi084,n305);
not gate_1813(n2027,n2026);
and gate_1814(n2028,pi046,n347);
and gate_1815(n2029,n304,n2028);
not gate_1816(n2030,n2029);
and gate_1817(n2031,n2027,n2030);
and gate_1818(n2032,n566,n2031);
and gate_1819(n2033,pi009,n346);
and gate_1820(n2034,n304,n2033);
and gate_1821(n2035,n324,n2034);
and gate_1822(n2036,n333,n2035);
not gate_1823(n2037,n2036);
and gate_1824(n2038,n351,n2037);
and gate_1825(n2039,n2032,n2038);
not gate_1826(n2040,n2039);
and gate_1827(n2041,n1506,n2040);
and gate_1828(n2042,n1507,n2041);
and gate_1829(n2043,n1451,n2042);
not gate_1830(n2044,n2043);
and gate_1831(n2045,n1452,n2040);
and gate_1832(n2046,n1508,n2045);
and gate_1833(n2047,pi005,n2046);
not gate_1834(n2048,n2047);
and gate_1835(n2049,n2044,n2048);
and gate_1836(n2050,n802,n1508);
and gate_1837(n2051,n245,n2050);
not gate_1838(n2052,n2051);
and gate_1839(n2053,n2049,n2052);
and gate_1840(n2054,n1509,n2040);
not gate_1841(n2055,n2054);
and gate_1842(n2056,n2053,n2055);
not gate_1843(po49,n2056);
and gate_1844(n2058,pi085,n305);
not gate_1845(n2059,n2058);
and gate_1846(n2060,pi047,n347);
and gate_1847(n2061,n304,n2060);
not gate_1848(n2062,n2061);
and gate_1849(n2063,n2059,n2062);
and gate_1850(n2064,n356,n2063);
and gate_1851(n2065,pi010,n346);
and gate_1852(n2066,n304,n2065);
and gate_1853(n2067,n324,n2066);
and gate_1854(n2068,n333,n2067);
not gate_1855(n2069,n2068);
and gate_1856(n2070,n351,n2069);
and gate_1857(n2071,n2064,n2070);
not gate_1858(n2072,n2071);
and gate_1859(n2073,n1506,n2072);
and gate_1860(n2074,n1507,n2073);
and gate_1861(n2075,n1451,n2074);
not gate_1862(n2076,n2075);
and gate_1863(n2077,n1452,n2072);
and gate_1864(n2078,n1508,n2077);
and gate_1865(n2079,pi005,n2078);
not gate_1866(n2080,n2079);
and gate_1867(n2081,n2076,n2080);
and gate_1868(n2082,n840,n1508);
and gate_1869(n2083,n245,n2082);
not gate_1870(n2084,n2083);
and gate_1871(n2085,n2081,n2084);
and gate_1872(n2086,n1509,n2072);
not gate_1873(n2087,n2086);
and gate_1874(n2088,n2085,n2087);
not gate_1875(po50,n2088);
and gate_1876(n2090,pi086,n305);
not gate_1877(n2091,n2090);
and gate_1878(n2092,pi048,n347);
and gate_1879(n2093,n304,n2092);
not gate_1880(n2094,n2093);
and gate_1881(n2095,n2091,n2094);
and gate_1882(n2096,n378,n2095);
and gate_1883(n2097,pi011,n346);
and gate_1884(n2098,n304,n2097);
and gate_1885(n2099,n324,n2098);
and gate_1886(n2100,n333,n2099);
not gate_1887(n2101,n2100);
and gate_1888(n2102,n351,n2101);
and gate_1889(n2103,n2096,n2102);
not gate_1890(n2104,n2103);
and gate_1891(n2105,n1506,n2104);
and gate_1892(n2106,n1507,n2105);
and gate_1893(n2107,n1451,n2106);
not gate_1894(n2108,n2107);
and gate_1895(n2109,n1452,n2104);
and gate_1896(n2110,n1508,n2109);
and gate_1897(n2111,pi005,n2110);
not gate_1898(n2112,n2111);
and gate_1899(n2113,n2108,n2112);
and gate_1900(n2114,n707,n1508);
and gate_1901(n2115,n245,n2114);
not gate_1902(n2116,n2115);
and gate_1903(n2117,n2113,n2116);
and gate_1904(n2118,n1509,n2104);
not gate_1905(n2119,n2118);
and gate_1906(n2120,n2117,n2119);
not gate_1907(po51,n2120);
and gate_1908(n2122,n325,n2002);
not gate_1909(n2123,n2122);
and gate_1910(n2124,pi041,n305);
not gate_1911(n2125,n2124);
and gate_1912(n2126,pi049,n347);
and gate_1913(n2127,n304,n2126);
not gate_1914(n2128,n2127);
and gate_1915(n2129,n2125,n2128);
and gate_1916(n2130,n2123,n2129);
and gate_1917(n2131,pi012,n346);
and gate_1918(n2132,n304,n2131);
and gate_1919(n2133,n324,n2132);
and gate_1920(n2134,n333,n2133);
not gate_1921(n2135,n2134);
and gate_1922(n2136,n351,n2135);
and gate_1923(n2137,n2130,n2136);
not gate_1924(n2138,n2137);
and gate_1925(n2139,n1506,n2138);
and gate_1926(n2140,n1507,n2139);
and gate_1927(n2141,n1451,n2140);
not gate_1928(n2142,n2141);
and gate_1929(n2143,n1452,n2138);
and gate_1930(n2144,n1508,n2143);
and gate_1931(n2145,pi005,n2144);
not gate_1932(n2146,n2145);
and gate_1933(n2147,n2142,n2146);
and gate_1934(n2148,n1452,n1508);
and gate_1935(n2149,n615,n2148);
not gate_1936(n2150,n2149);
and gate_1937(n2151,n2147,n2150);
and gate_1938(n2152,n1509,n2138);
not gate_1939(n2153,n2152);
and gate_1940(n2154,n2151,n2153);
not gate_1941(po52,n2154);
and gate_1942(n2156,n325,n2034);
not gate_1943(n2157,n2156);
and gate_1944(n2158,pi042,n305);
not gate_1945(n2159,n2158);
and gate_1946(n2160,pi050,n347);
and gate_1947(n2161,n304,n2160);
not gate_1948(n2162,n2161);
and gate_1949(n2163,n2159,n2162);
and gate_1950(n2164,n2157,n2163);
and gate_1951(n2165,pi013,n346);
and gate_1952(n2166,n304,n2165);
and gate_1953(n2167,n324,n2166);
and gate_1954(n2168,n333,n2167);
not gate_1955(n2169,n2168);
and gate_1956(n2170,n351,n2169);
and gate_1957(n2171,n2164,n2170);
not gate_1958(n2172,n2171);
and gate_1959(n2173,n1509,n2172);
not gate_1960(n2174,n2173);
and gate_1961(n2175,n1506,n2172);
and gate_1962(n2176,n1507,n2175);
and gate_1963(n2177,n1451,n2176);
not gate_1964(n2178,n2177);
and gate_1965(n2179,pi005,n2172);
not gate_1966(n2180,n2179);
and gate_1967(n2181,n643,n2180);
not gate_1968(n2182,n2181);
and gate_1969(n2183,n2148,n2182);
not gate_1970(n2184,n2183);
and gate_1971(n2185,n2178,n2184);
and gate_1972(n2186,n2174,n2185);
not gate_1973(po53,n2186);
and gate_1974(n2188,n325,n2066);
not gate_1975(n2189,n2188);
and gate_1976(n2190,pi043,n305);
not gate_1977(n2191,n2190);
and gate_1978(n2192,pi051,n347);
and gate_1979(n2193,n304,n2192);
not gate_1980(n2194,n2193);
and gate_1981(n2195,n2191,n2194);
and gate_1982(n2196,n2189,n2195);
and gate_1983(n2197,pi014,n346);
and gate_1984(n2198,n304,n2197);
and gate_1985(n2199,n324,n2198);
and gate_1986(n2200,n333,n2199);
not gate_1987(n2201,n2200);
and gate_1988(n2202,n351,n2201);
and gate_1989(n2203,n2196,n2202);
not gate_1990(n2204,n2203);
and gate_1991(n2205,n1509,n2204);
not gate_1992(n2206,n2205);
and gate_1993(n2207,n1506,n2204);
and gate_1994(n2208,n1507,n2207);
and gate_1995(n2209,n1451,n2208);
not gate_1996(n2210,n2209);
and gate_1997(n2211,pi005,n2204);
not gate_1998(n2212,n2211);
and gate_1999(n2213,n610,n2212);
not gate_2000(n2214,n2213);
and gate_2001(n2215,n2148,n2214);
not gate_2002(n2216,n2215);
and gate_2003(n2217,n2210,n2216);
and gate_2004(n2218,n2206,n2217);
not gate_2005(po54,n2218);
and gate_2006(n2220,n325,n2098);
not gate_2007(n2221,n2220);
and gate_2008(n2222,pi044,n305);
not gate_2009(n2223,n2222);
and gate_2010(n2224,pi087,n347);
and gate_2011(n2225,n304,n2224);
not gate_2012(n2226,n2225);
and gate_2013(n2227,n2223,n2226);
and gate_2014(n2228,n2221,n2227);
and gate_2015(n2229,pi015,n346);
and gate_2016(n2230,n304,n2229);
and gate_2017(n2231,n324,n2230);
and gate_2018(n2232,n333,n2231);
not gate_2019(n2233,n2232);
and gate_2020(n2234,n351,n2233);
and gate_2021(n2235,n2228,n2234);
not gate_2022(n2236,n2235);
and gate_2023(n2237,n1506,n2236);
and gate_2024(n2238,n1507,n2237);
and gate_2025(n2239,n1451,n2238);
not gate_2026(n2240,n2239);
and gate_2027(n2241,pi005,n2236);
and gate_2028(n2242,n2148,n2241);
not gate_2029(n2243,n2242);
and gate_2030(n2244,n2240,n2243);
and gate_2031(n2245,n447,n2148);
and gate_2032(n2246,n245,n2245);
not gate_2033(n2247,n2246);
and gate_2034(n2248,n2244,n2247);
and gate_2035(n2249,n1509,n2236);
not gate_2036(n2250,n2249);
and gate_2037(n2251,n2248,n2250);
not gate_2038(po55,n2251);
and gate_2039(n2253,n325,n2132);
not gate_2040(n2254,n2253);
and gate_2041(n2255,pi045,n305);
not gate_2042(n2256,n2255);
and gate_2043(n2257,pi009,n347);
and gate_2044(n2258,n304,n2257);
not gate_2045(n2259,n2258);
and gate_2046(n2260,n2256,n2259);
and gate_2047(n2261,n2254,n2260);
and gate_2048(n2262,pi016,n346);
and gate_2049(n2263,n304,n2262);
and gate_2050(n2264,n324,n2263);
and gate_2051(n2265,n333,n2264);
not gate_2052(n2266,n2265);
and gate_2053(n2267,n351,n2266);
and gate_2054(n2268,n2261,n2267);
not gate_2055(n2269,n2268);
and gate_2056(n2270,n1506,n2269);
and gate_2057(n2271,n1507,n2270);
and gate_2058(n2272,n1451,n2271);
not gate_2059(n2273,n2272);
and gate_2060(n2274,pi005,n2269);
and gate_2061(n2275,n2148,n2274);
not gate_2062(n2276,n2275);
and gate_2063(n2277,n2273,n2276);
and gate_2064(n2278,n458,n2148);
and gate_2065(n2279,n245,n2278);
not gate_2066(n2280,n2279);
and gate_2067(n2281,n2277,n2280);
and gate_2068(n2282,n1509,n2269);
not gate_2069(n2283,n2282);
and gate_2070(n2284,n2281,n2283);
not gate_2071(po56,n2284);
and gate_2072(n2286,n325,n2166);
not gate_2073(n2287,n2286);
and gate_2074(n2288,pi046,n305);
not gate_2075(n2289,n2288);
and gate_2076(n2290,pi010,n347);
and gate_2077(n2291,n304,n2290);
not gate_2078(n2292,n2291);
and gate_2079(n2293,n2289,n2292);
and gate_2080(n2294,n2287,n2293);
and gate_2081(n2295,pi017,n346);
and gate_2082(n2296,n304,n2295);
and gate_2083(n2297,n324,n2296);
and gate_2084(n2298,n333,n2297);
not gate_2085(n2299,n2298);
and gate_2086(n2300,n351,n2299);
and gate_2087(n2301,n2294,n2300);
not gate_2088(n2302,n2301);
and gate_2089(n2303,n1509,n2302);
not gate_2090(n2304,n2303);
and gate_2091(n2305,n1506,n2302);
and gate_2092(n2306,n1507,n2305);
and gate_2093(n2307,n1451,n2306);
not gate_2094(n2308,n2307);
and gate_2095(n2309,pi005,n2302);
not gate_2096(n2310,n2309);
and gate_2097(n2311,n485,n2310);
not gate_2098(n2312,n2311);
and gate_2099(n2313,n2148,n2312);
not gate_2100(n2314,n2313);
and gate_2101(n2315,n2308,n2314);
and gate_2102(n2316,n2304,n2315);
not gate_2103(po57,n2316);
and gate_2104(n2318,n325,n2198);
not gate_2105(n2319,n2318);
and gate_2106(n2320,pi047,n305);
not gate_2107(n2321,n2320);
and gate_2108(n2322,pi011,n347);
and gate_2109(n2323,n304,n2322);
not gate_2110(n2324,n2323);
and gate_2111(n2325,n2321,n2324);
and gate_2112(n2326,n2319,n2325);
and gate_2113(n2327,pi018,n346);
and gate_2114(n2328,n304,n2327);
and gate_2115(n2329,n324,n2328);
and gate_2116(n2330,n333,n2329);
not gate_2117(n2331,n2330);
and gate_2118(n2332,n351,n2331);
and gate_2119(n2333,n2326,n2332);
not gate_2120(n2334,n2333);
and gate_2121(n2335,n1509,n2334);
not gate_2122(n2336,n2335);
and gate_2123(n2337,n1506,n2334);
and gate_2124(n2338,n1507,n2337);
and gate_2125(n2339,n1451,n2338);
not gate_2126(n2340,n2339);
and gate_2127(n2341,pi005,n2334);
not gate_2128(n2342,n2341);
and gate_2129(n2343,n509,n2342);
not gate_2130(n2344,n2343);
and gate_2131(n2345,n2148,n2344);
not gate_2132(n2346,n2345);
and gate_2133(n2347,n2340,n2346);
and gate_2134(n2348,n2336,n2347);
not gate_2135(po58,n2348);
and gate_2136(n2350,n325,n2230);
not gate_2137(n2351,n2350);
and gate_2138(n2352,pi048,n305);
not gate_2139(n2353,n2352);
and gate_2140(n2354,pi012,n347);
and gate_2141(n2355,n304,n2354);
not gate_2142(n2356,n2355);
and gate_2143(n2357,n2353,n2356);
and gate_2144(n2358,n2351,n2357);
and gate_2145(n2359,pi019,n346);
and gate_2146(n2360,n304,n2359);
and gate_2147(n2361,n324,n2360);
and gate_2148(n2362,n333,n2361);
not gate_2149(n2363,n2362);
and gate_2150(n2364,n351,n2363);
and gate_2151(n2365,n2358,n2364);
not gate_2152(n2366,n2365);
and gate_2153(n2367,n1509,n2366);
not gate_2154(n2368,n2367);
and gate_2155(n2369,n1506,n2366);
and gate_2156(n2370,n1507,n2369);
and gate_2157(n2371,n1451,n2370);
not gate_2158(n2372,n2371);
and gate_2159(n2373,pi005,n2366);
not gate_2160(n2374,n2373);
and gate_2161(n2375,n533,n2374);
not gate_2162(n2376,n2375);
and gate_2163(n2377,n2148,n2376);
not gate_2164(n2378,n2377);
and gate_2165(n2379,n2372,n2378);
and gate_2166(n2380,n2368,n2379);
not gate_2167(po59,n2380);
and gate_2168(n2382,n325,n2263);
not gate_2169(n2383,n2382);
and gate_2170(n2384,pi049,n305);
not gate_2171(n2385,n2384);
and gate_2172(n2386,pi013,n347);
and gate_2173(n2387,n304,n2386);
not gate_2174(n2388,n2387);
and gate_2175(n2389,n2385,n2388);
and gate_2176(n2390,n2383,n2389);
and gate_2177(n2391,n324,n912);
and gate_2178(n2392,n333,n2391);
not gate_2179(n2393,n2392);
and gate_2180(n2394,n351,n2393);
and gate_2181(n2395,n2390,n2394);
not gate_2182(n2396,n2395);
and gate_2183(n2397,n1509,n2396);
not gate_2184(n2398,n2397);
and gate_2185(n2399,n1506,n2396);
and gate_2186(n2400,n1507,n2399);
and gate_2187(n2401,n1451,n2400);
not gate_2188(n2402,n2401);
and gate_2189(n2403,pi005,n2396);
not gate_2190(n2404,n2403);
and gate_2191(n2405,n557,n2404);
not gate_2192(n2406,n2405);
and gate_2193(n2407,n2148,n2406);
not gate_2194(n2408,n2407);
and gate_2195(n2409,n2402,n2408);
and gate_2196(n2410,n2398,n2409);
not gate_2197(po60,n2410);
and gate_2198(n2412,n325,n2296);
not gate_2199(n2413,n2412);
and gate_2200(n2414,pi050,n305);
not gate_2201(n2415,n2414);
and gate_2202(n2416,pi014,n347);
and gate_2203(n2417,n304,n2416);
not gate_2204(n2418,n2417);
and gate_2205(n2419,n2415,n2418);
and gate_2206(n2420,n2413,n2419);
and gate_2207(n2421,n324,n950);
and gate_2208(n2422,n333,n2421);
not gate_2209(n2423,n2422);
and gate_2210(n2424,n351,n2423);
and gate_2211(n2425,n2420,n2424);
not gate_2212(n2426,n2425);
and gate_2213(n2427,n1506,n2426);
and gate_2214(n2428,n1507,n2427);
and gate_2215(n2429,n1451,n2428);
not gate_2216(n2430,n2429);
and gate_2217(n2431,pi005,n2426);
and gate_2218(n2432,n2148,n2431);
not gate_2219(n2433,n2432);
and gate_2220(n2434,n2430,n2433);
and gate_2221(n2435,pi094,n2148);
and gate_2222(n2436,n245,n2435);
not gate_2223(n2437,n2436);
and gate_2224(n2438,n2434,n2437);
and gate_2225(n2439,n1509,n2426);
not gate_2226(n2440,n2439);
and gate_2227(n2441,n2438,n2440);
not gate_2228(po61,n2441);
and gate_2229(n2443,n325,n2328);
not gate_2230(n2444,n2443);
and gate_2231(n2445,pi051,n305);
not gate_2232(n2446,n2445);
and gate_2233(n2447,pi015,n347);
and gate_2234(n2448,n304,n2447);
not gate_2235(n2449,n2448);
and gate_2236(n2450,n2446,n2449);
and gate_2237(n2451,n2444,n2450);
and gate_2238(n2452,n324,n988);
and gate_2239(n2453,n333,n2452);
not gate_2240(n2454,n2453);
and gate_2241(n2455,n351,n2454);
and gate_2242(n2456,n2451,n2455);
not gate_2243(n2457,n2456);
and gate_2244(n2458,n1506,n2457);
and gate_2245(n2459,n1507,n2458);
and gate_2246(n2460,n1451,n2459);
not gate_2247(n2461,n2460);
and gate_2248(n2462,pi005,n2457);
and gate_2249(n2463,n2148,n2462);
not gate_2250(n2464,n2463);
and gate_2251(n2465,n2461,n2464);
and gate_2252(n2466,pi096,n2148);
and gate_2253(n2467,n245,n2466);
not gate_2254(n2468,n2467);
and gate_2255(n2469,n2465,n2468);
and gate_2256(n2470,n1509,n2457);
not gate_2257(n2471,n2470);
and gate_2258(n2472,n2469,n2471);
not gate_2259(po62,n2472);
and gate_2260(n2474,n325,n2360);
not gate_2261(n2475,n2474);
and gate_2262(n2476,pi087,n305);
not gate_2263(n2477,n2476);
and gate_2264(n2478,pi016,n347);
and gate_2265(n2479,n304,n2478);
not gate_2266(n2480,n2479);
and gate_2267(n2481,n2477,n2480);
and gate_2268(n2482,n2475,n2481);
and gate_2269(n2483,n324,n1026);
and gate_2270(n2484,n333,n2483);
not gate_2271(n2485,n2484);
and gate_2272(n2486,n351,n2485);
and gate_2273(n2487,n2482,n2486);
not gate_2274(n2488,n2487);
and gate_2275(n2489,n1506,n2488);
and gate_2276(n2490,n1507,n2489);
and gate_2277(n2491,n1451,n2490);
not gate_2278(n2492,n2491);
and gate_2279(n2493,pi005,n2488);
and gate_2280(n2494,n2148,n2493);
not gate_2281(n2495,n2494);
and gate_2282(n2496,n2492,n2495);
and gate_2283(n2497,pi090,n2148);
and gate_2284(n2498,n245,n2497);
not gate_2285(n2499,n2498);
and gate_2286(n2500,n2496,n2499);
and gate_2287(n2501,n1509,n2488);
not gate_2288(n2502,n2501);
and gate_2289(n2503,n2500,n2502);
not gate_2290(po63,n2503);
and gate_2291(n2505,n215,n226);
and gate_2292(n2506,n216,n2505);
and gate_2293(n2507,n225,n2506);
and gate_2294(n2508,n227,n2507);
and gate_2295(n2509,n342,n2508);
not gate_2296(n2510,n2509);
and gate_2297(n2511,n220,n854);
and gate_2298(n2512,n218,n2511);
not gate_2299(n2513,n2512);
and gate_2300(n2514,pi007,n853);
not gate_2301(n2515,n2514);
and gate_2302(n2516,pi108,n2510);
and gate_2303(n2517,n2515,n2516);
and gate_2304(n2518,n2513,n2517);
and gate_2305(n2519,n245,n2518);
not gate_2306(n2520,n2519);
and gate_2307(n2521,n2510,n2520);
and gate_2308(n2522,n219,n2515);
and gate_2309(n2523,n2513,n2522);
not gate_2310(n2524,n2523);
and gate_2311(n2525,pi067,n2524);
not gate_2312(n2526,n2525);
and gate_2313(n2527,n2521,n2526);
not gate_2314(po64,n2527);
and gate_2315(n2529,pi068,n2524);
not gate_2316(n2530,n2529);
and gate_2317(n2531,pi109,n245);
and gate_2318(n2532,n2523,n2531);
not gate_2319(n2533,n2532);
and gate_2320(n2534,n2510,n2533);
and gate_2321(n2535,n2530,n2534);
not gate_2322(po65,n2535);
and gate_2323(n2537,pi069,n2524);
not gate_2324(n2538,n2537);
and gate_2325(n2539,pi106,n245);
and gate_2326(n2540,n2523,n2539);
not gate_2327(n2541,n2540);
and gate_2328(n2542,n2510,n2541);
and gate_2329(n2543,n2538,n2542);
not gate_2330(po66,n2543);
and gate_2331(n2545,pi070,n2524);
not gate_2332(n2546,n2545);
and gate_2333(n2547,pi104,n245);
and gate_2334(n2548,n2523,n2547);
not gate_2335(n2549,n2548);
and gate_2336(n2550,n2510,n2549);
and gate_2337(n2551,n2546,n2550);
not gate_2338(po67,n2551);
and gate_2339(n2553,pi071,n2524);
not gate_2340(n2554,n2553);
and gate_2341(n2555,pi105,n245);
and gate_2342(n2556,n2523,n2555);
not gate_2343(n2557,n2556);
and gate_2344(n2558,n2510,n2557);
and gate_2345(n2559,n2554,n2558);
not gate_2346(po68,n2559);
and gate_2347(n2561,pi072,n2524);
not gate_2348(n2562,n2561);
and gate_2349(n2563,pi103,n245);
and gate_2350(n2564,n2523,n2563);
not gate_2351(n2565,n2564);
and gate_2352(n2566,n2510,n2565);
and gate_2353(n2567,n2562,n2566);
not gate_2354(po69,n2567);
and gate_2355(n2569,pi073,n2524);
not gate_2356(n2570,n2569);
and gate_2357(n2571,pi097,n245);
and gate_2358(n2572,n2523,n2571);
not gate_2359(n2573,n2572);
and gate_2360(n2574,n2510,n2573);
and gate_2361(n2575,n2570,n2574);
not gate_2362(po70,n2575);
and gate_2363(n2577,pi074,n2524);
not gate_2364(n2578,n2577);
and gate_2365(n2579,pi098,n245);
and gate_2366(n2580,n2523,n2579);
not gate_2367(n2581,n2580);
and gate_2368(n2582,n2510,n2581);
and gate_2369(n2583,n2578,n2582);
not gate_2370(po71,n2583);
and gate_2371(n2585,pi075,n2524);
not gate_2372(n2586,n2585);
and gate_2373(n2587,pi099,n245);
and gate_2374(n2588,n2523,n2587);
not gate_2375(n2589,n2588);
and gate_2376(n2590,n2510,n2589);
and gate_2377(n2591,n2586,n2590);
not gate_2378(po72,n2591);
and gate_2379(n2593,pi076,n2524);
not gate_2380(n2594,n2593);
and gate_2381(n2595,pi100,n245);
and gate_2382(n2596,n2523,n2595);
not gate_2383(n2597,n2596);
and gate_2384(n2598,n2510,n2597);
and gate_2385(n2599,n2594,n2598);
not gate_2386(po73,n2599);
and gate_2387(n2601,pi077,n2524);
not gate_2388(n2602,n2601);
and gate_2389(n2603,pi101,n245);
and gate_2390(n2604,n2523,n2603);
not gate_2391(n2605,n2604);
and gate_2392(n2606,n2510,n2605);
and gate_2393(n2607,n2602,n2606);
not gate_2394(po74,n2607);
and gate_2395(n2609,pi078,n2524);
not gate_2396(n2610,n2609);
and gate_2397(n2611,pi102,n245);
and gate_2398(n2612,n2523,n2611);
not gate_2399(n2613,n2612);
and gate_2400(n2614,n2510,n2613);
and gate_2401(n2615,n2610,n2614);
not gate_2402(po75,n2615);
and gate_2403(n2617,pi079,n2524);
not gate_2404(n2618,n2617);
and gate_2405(n2619,pi094,n245);
and gate_2406(n2620,n2523,n2619);
not gate_2407(n2621,n2620);
and gate_2408(n2622,n2510,n2621);
and gate_2409(n2623,n2618,n2622);
not gate_2410(po76,n2623);
and gate_2411(n2625,pi080,n2524);
not gate_2412(n2626,n2625);
and gate_2413(n2627,pi096,n245);
and gate_2414(n2628,n2523,n2627);
not gate_2415(n2629,n2628);
and gate_2416(n2630,n2510,n2629);
and gate_2417(n2631,n2626,n2630);
not gate_2418(po77,n2631);
and gate_2419(n2633,pi081,n2524);
not gate_2420(n2634,n2633);
and gate_2421(n2635,pi090,n245);
and gate_2422(n2636,n2523,n2635);
not gate_2423(n2637,n2636);
and gate_2424(n2638,n2510,n2637);
and gate_2425(n2639,n2634,n2638);
not gate_2426(po78,n2639);
and gate_2427(n2641,n278,n320);
and gate_2428(n2642,n269,n2641);
not gate_2429(n2643,n2642);
and gate_2430(n2644,pi007,n227);
not gate_2431(n2645,n2644);
and gate_2432(n2646,n222,n2644);
not gate_2433(n2647,n2646);
and gate_2434(n2648,pi126,n2646);
not gate_2435(n2649,n2648);
and gate_2436(n2650,n246,n280);
and gate_2437(n2651,n2647,n2650);
and gate_2438(n2652,n320,n2651);
and gate_2439(n2653,n269,n2652);
not gate_2440(n2654,n2653);
and gate_2441(n2655,n2649,n2654);
and gate_2442(n2656,n2643,n2655);
and gate_2443(n2657,n268,n320);
not gate_2444(n2658,n2657);
and gate_2445(n2659,pi127,n320);
and gate_2446(n2660,pi005,n2659);
and gate_2447(n2661,n2647,n2660);
not gate_2448(n2662,n2661);
and gate_2449(n2663,n2658,n2662);
and gate_2450(n2664,n2656,n2663);
not gate_2451(po79,n2664);
and gate_2452(n2666,pi128,n2644);
not gate_2453(n2667,n2666);
and gate_2454(n2668,n223,n319);
not gate_2455(n2669,n2668);
and gate_2456(n2670,n2645,n2668);
not gate_2457(n2671,n2670);
and gate_2458(n2672,n2667,n2671);
and gate_2459(n2673,pi129,n2669);
and gate_2460(n2674,pi005,n2673);
not gate_2461(n2675,n2674);
and gate_2462(n2676,n2672,n2675);
not gate_2463(po80,n2676);
endmodule
