// Verilog File 
module c1355 (G1gat,G8gat,G15gat,G22gat,G29gat,G36gat,G43gat,G50gat,G57gat,
G64gat,G71gat,G78gat,G85gat,G92gat,G99gat,G106gat,G113gat,G120gat,G127gat,
G134gat,G141gat,G148gat,G155gat,G162gat,G169gat,G176gat,G183gat,G190gat,G197gat,
G204gat,G211gat,G218gat,G225gat,G226gat,G227gat,G228gat,G229gat,G230gat,G231gat,
G232gat,G233gat,G1324gat,G1325gat,G1326gat,G1327gat,G1328gat,G1329gat,G1330gat,G1331gat,
G1332gat,G1333gat,G1334gat,G1335gat,G1336gat,G1337gat,G1338gat,G1339gat,G1340gat,G1341gat,
G1342gat,G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,
G1352gat,G1353gat,G1354gat,G1355gat);

input G1gat,G8gat,G15gat,G22gat,G29gat,G36gat,G43gat,G50gat,G57gat,
G64gat,G71gat,G78gat,G85gat,G92gat,G99gat,G106gat,G113gat,G120gat,G127gat,
G134gat,G141gat,G148gat,G155gat,G162gat,G169gat,G176gat,G183gat,G190gat,G197gat,
G204gat,G211gat,G218gat,G225gat,G226gat,G227gat,G228gat,G229gat,G230gat,G231gat,
G232gat,G233gat;

output G1324gat,G1325gat,G1326gat,G1327gat,G1328gat,G1329gat,G1330gat,G1331gat,G1332gat,
G1333gat,G1334gat,G1335gat,G1336gat,G1337gat,G1338gat,G1339gat,G1340gat,G1341gat,G1342gat,
G1343gat,G1344gat,G1345gat,G1346gat,G1347gat,G1348gat,G1349gat,G1350gat,G1351gat,G1352gat,
G1353gat,G1354gat,G1355gat;

wire G242gat,G245gat,G248gat,G251gat,G254gat,G257gat,G260gat,G263gat,G266gat,
G269gat,G272gat,G275gat,G278gat,G281gat,G284gat,G287gat,G290gat,G293gat,G296gat,
G299gat,G302gat,G305gat,G308gat,G311gat,G314gat,G317gat,G320gat,G323gat,G326gat,
G329gat,G332gat,G335gat,G338gat,G341gat,G344gat,G347gat,G350gat,G353gat,G356gat,
G359gat,G362gat,G363gat,G364gat,G365gat,G366gat,G367gat,G368gat,G369gat,G370gat,
G371gat,G372gat,G373gat,G374gat,G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,
G381gat,G382gat,G383gat,G384gat,G385gat,G386gat,G387gat,G388gat,G389gat,G390gat,
G391gat,G392gat,G393gat,G394gat,G395gat,G396gat,G397gat,G398gat,G399gat,G400gat,
G401gat,G402gat,G403gat,G404gat,G405gat,G406gat,G407gat,G408gat,G409gat,G410gat,
G411gat,G412gat,G413gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,
G421gat,G422gat,G423gat,G424gat,G425gat,G426gat,G429gat,G432gat,G435gat,G438gat,
G441gat,G444gat,G447gat,G450gat,G453gat,G456gat,G459gat,G462gat,G465gat,G468gat,
G471gat,G474gat,G477gat,G480gat,G483gat,G486gat,G489gat,G492gat,G495gat,G498gat,
G501gat,G504gat,G507gat,G510gat,G513gat,G516gat,G519gat,G522gat,G525gat,G528gat,
G531gat,G534gat,G537gat,G540gat,G543gat,G546gat,G549gat,G552gat,G555gat,G558gat,
G561gat,G564gat,G567gat,G570gat,G571gat,G572gat,G573gat,G574gat,G575gat,G576gat,
G577gat,G578gat,G579gat,G580gat,G581gat,G582gat,G583gat,G584gat,G585gat,G586gat,
G587gat,G588gat,G589gat,G590gat,G591gat,G592gat,G593gat,G594gat,G595gat,G596gat,
G597gat,G598gat,G599gat,G600gat,G601gat,G602gat,G607gat,G612gat,G617gat,G622gat,
G627gat,G632gat,G637gat,G642gat,G645gat,G648gat,G651gat,G654gat,G657gat,G660gat,
G663gat,G666gat,G669gat,G672gat,G675gat,G678gat,G681gat,G684gat,G687gat,G690gat,
G691gat,G692gat,G693gat,G694gat,G695gat,G696gat,G697gat,G698gat,G699gat,G700gat,
G701gat,G702gat,G703gat,G704gat,G705gat,G706gat,G709gat,G712gat,G715gat,G718gat,
G721gat,G724gat,G727gat,G730gat,G733gat,G736gat,G739gat,G742gat,G745gat,G748gat,
G751gat,G754gat,G755gat,G756gat,G757gat,G758gat,G759gat,G760gat,G761gat,G762gat,
G763gat,G764gat,G765gat,G766gat,G767gat,G768gat,G769gat,G770gat,G773gat,G776gat,
G779gat,G782gat,G785gat,G788gat,G791gat,G794gat,G797gat,G800gat,G803gat,G806gat,
G809gat,G812gat,G815gat,G818gat,G819gat,G820gat,G821gat,G822gat,G823gat,G824gat,
G825gat,G826gat,G827gat,G828gat,G829gat,G830gat,G831gat,G832gat,G833gat,G834gat,
G847gat,G860gat,G873gat,G886gat,G899gat,G912gat,G925gat,G938gat,G939gat,G940gat,
G941gat,G942gat,G943gat,G944gat,G945gat,G946gat,G947gat,G948gat,G949gat,G950gat,
G951gat,G952gat,G953gat,G954gat,G955gat,G956gat,G957gat,G958gat,G959gat,G960gat,
G961gat,G962gat,G963gat,G964gat,G965gat,G966gat,G967gat,G968gat,G969gat,G970gat,
G971gat,G972gat,G973gat,G974gat,G975gat,G976gat,G977gat,G978gat,G979gat,G980gat,
G981gat,G982gat,G983gat,G984gat,G985gat,G986gat,G991gat,G996gat,G1001gat,G1006gat,
G1011gat,G1016gat,G1021gat,G1026gat,G1031gat,G1036gat,G1039gat,G1042gat,G1045gat,G1048gat,
G1051gat,G1054gat,G1057gat,G1060gat,G1063gat,G1066gat,G1069gat,G1072gat,G1075gat,G1078gat,
G1081gat,G1084gat,G1087gat,G1090gat,G1093gat,G1096gat,G1099gat,G1102gat,G1105gat,G1108gat,
G1111gat,G1114gat,G1117gat,G1120gat,G1123gat,G1126gat,G1129gat,G1132gat,G1135gat,G1138gat,
G1141gat,G1144gat,G1147gat,G1150gat,G1153gat,G1156gat,G1159gat,G1162gat,G1165gat,G1168gat,
G1171gat,G1174gat,G1177gat,G1180gat,G1183gat,G1186gat,G1189gat,G1192gat,G1195gat,G1198gat,
G1201gat,G1204gat,G1207gat,G1210gat,G1213gat,G1216gat,G1219gat,G1222gat,G1225gat,G1228gat,
G1229gat,G1230gat,G1231gat,G1232gat,G1233gat,G1234gat,G1235gat,G1236gat,G1237gat,G1238gat,
G1239gat,G1240gat,G1241gat,G1242gat,G1243gat,G1244gat,G1245gat,G1246gat,G1247gat,G1248gat,
G1249gat,G1250gat,G1251gat,G1252gat,G1253gat,G1254gat,G1255gat,G1256gat,G1257gat,G1258gat,
G1259gat,G1260gat,G1261gat,G1262gat,G1263gat,G1264gat,G1265gat,G1266gat,G1267gat,G1268gat,
G1269gat,G1270gat,G1271gat,G1272gat,G1273gat,G1274gat,G1275gat,G1276gat,G1277gat,G1278gat,
G1279gat,G1280gat,G1281gat,G1282gat,G1283gat,G1284gat,G1285gat,G1286gat,G1287gat,G1288gat,
G1289gat,G1290gat,G1291gat,G1292gat,G1293gat,G1294gat,G1295gat,G1296gat,G1297gat,G1298gat,
G1299gat,G1300gat,G1301gat,G1302gat,G1303gat,G1304gat,G1305gat,G1306gat,G1307gat,G1308gat,
G1309gat,G1310gat,G1311gat,G1312gat,G1313gat,G1314gat,G1315gat,G1316gat,G1317gat,G1318gat,
G1319gat,G1320gat,G1321gat,G1322gat,G1323gat;
and gate_0(G242gat,G225gat,G233gat);
and gate_1(G245gat,G226gat,G233gat);
and gate_2(G248gat,G227gat,G233gat);
and gate_3(G251gat,G228gat,G233gat);
and gate_4(G254gat,G229gat,G233gat);
and gate_5(G257gat,G230gat,G233gat);
and gate_6(G260gat,G231gat,G233gat);
and gate_7(G263gat,G232gat,G233gat);
nand gate_8(G266gat,G1gat,G8gat);
nand gate_9(G269gat,G15gat,G22gat);
nand gate_10(G272gat,G29gat,G36gat);
nand gate_11(G275gat,G43gat,G50gat);
nand gate_12(G278gat,G57gat,G64gat);
nand gate_13(G281gat,G71gat,G78gat);
nand gate_14(G284gat,G85gat,G92gat);
nand gate_15(G287gat,G99gat,G106gat);
nand gate_16(G290gat,G113gat,G120gat);
nand gate_17(G293gat,G127gat,G134gat);
nand gate_18(G296gat,G141gat,G148gat);
nand gate_19(G299gat,G155gat,G162gat);
nand gate_20(G302gat,G169gat,G176gat);
nand gate_21(G305gat,G183gat,G190gat);
nand gate_22(G308gat,G197gat,G204gat);
nand gate_23(G311gat,G211gat,G218gat);
nand gate_24(G314gat,G1gat,G29gat);
nand gate_25(G317gat,G57gat,G85gat);
nand gate_26(G320gat,G8gat,G36gat);
nand gate_27(G323gat,G64gat,G92gat);
nand gate_28(G326gat,G15gat,G43gat);
nand gate_29(G329gat,G71gat,G99gat);
nand gate_30(G332gat,G22gat,G50gat);
nand gate_31(G335gat,G78gat,G106gat);
nand gate_32(G338gat,G113gat,G141gat);
nand gate_33(G341gat,G169gat,G197gat);
nand gate_34(G344gat,G120gat,G148gat);
nand gate_35(G347gat,G176gat,G204gat);
nand gate_36(G350gat,G127gat,G155gat);
nand gate_37(G353gat,G183gat,G211gat);
nand gate_38(G356gat,G134gat,G162gat);
nand gate_39(G359gat,G190gat,G218gat);
nand gate_40(G362gat,G1gat,G266gat);
nand gate_41(G363gat,G8gat,G266gat);
nand gate_42(G364gat,G15gat,G269gat);
nand gate_43(G365gat,G22gat,G269gat);
nand gate_44(G366gat,G29gat,G272gat);
nand gate_45(G367gat,G36gat,G272gat);
nand gate_46(G368gat,G43gat,G275gat);
nand gate_47(G369gat,G50gat,G275gat);
nand gate_48(G370gat,G57gat,G278gat);
nand gate_49(G371gat,G64gat,G278gat);
nand gate_50(G372gat,G71gat,G281gat);
nand gate_51(G373gat,G78gat,G281gat);
nand gate_52(G374gat,G85gat,G284gat);
nand gate_53(G375gat,G92gat,G284gat);
nand gate_54(G376gat,G99gat,G287gat);
nand gate_55(G377gat,G106gat,G287gat);
nand gate_56(G378gat,G113gat,G290gat);
nand gate_57(G379gat,G120gat,G290gat);
nand gate_58(G380gat,G127gat,G293gat);
nand gate_59(G381gat,G134gat,G293gat);
nand gate_60(G382gat,G141gat,G296gat);
nand gate_61(G383gat,G148gat,G296gat);
nand gate_62(G384gat,G155gat,G299gat);
nand gate_63(G385gat,G162gat,G299gat);
nand gate_64(G386gat,G169gat,G302gat);
nand gate_65(G387gat,G176gat,G302gat);
nand gate_66(G388gat,G183gat,G305gat);
nand gate_67(G389gat,G190gat,G305gat);
nand gate_68(G390gat,G197gat,G308gat);
nand gate_69(G391gat,G204gat,G308gat);
nand gate_70(G392gat,G211gat,G311gat);
nand gate_71(G393gat,G218gat,G311gat);
nand gate_72(G394gat,G1gat,G314gat);
nand gate_73(G395gat,G29gat,G314gat);
nand gate_74(G396gat,G57gat,G317gat);
nand gate_75(G397gat,G85gat,G317gat);
nand gate_76(G398gat,G8gat,G320gat);
nand gate_77(G399gat,G36gat,G320gat);
nand gate_78(G400gat,G64gat,G323gat);
nand gate_79(G401gat,G92gat,G323gat);
nand gate_80(G402gat,G15gat,G326gat);
nand gate_81(G403gat,G43gat,G326gat);
nand gate_82(G404gat,G71gat,G329gat);
nand gate_83(G405gat,G99gat,G329gat);
nand gate_84(G406gat,G22gat,G332gat);
nand gate_85(G407gat,G50gat,G332gat);
nand gate_86(G408gat,G78gat,G335gat);
nand gate_87(G409gat,G106gat,G335gat);
nand gate_88(G410gat,G113gat,G338gat);
nand gate_89(G411gat,G141gat,G338gat);
nand gate_90(G412gat,G169gat,G341gat);
nand gate_91(G413gat,G197gat,G341gat);
nand gate_92(G414gat,G120gat,G344gat);
nand gate_93(G415gat,G148gat,G344gat);
nand gate_94(G416gat,G176gat,G347gat);
nand gate_95(G417gat,G204gat,G347gat);
nand gate_96(G418gat,G127gat,G350gat);
nand gate_97(G419gat,G155gat,G350gat);
nand gate_98(G420gat,G183gat,G353gat);
nand gate_99(G421gat,G211gat,G353gat);
nand gate_100(G422gat,G134gat,G356gat);
nand gate_101(G423gat,G162gat,G356gat);
nand gate_102(G424gat,G190gat,G359gat);
nand gate_103(G425gat,G218gat,G359gat);
nand gate_104(G426gat,G362gat,G363gat);
nand gate_105(G429gat,G364gat,G365gat);
nand gate_106(G432gat,G366gat,G367gat);
nand gate_107(G435gat,G368gat,G369gat);
nand gate_108(G438gat,G370gat,G371gat);
nand gate_109(G441gat,G372gat,G373gat);
nand gate_110(G444gat,G374gat,G375gat);
nand gate_111(G447gat,G376gat,G377gat);
nand gate_112(G450gat,G378gat,G379gat);
nand gate_113(G453gat,G380gat,G381gat);
nand gate_114(G456gat,G382gat,G383gat);
nand gate_115(G459gat,G384gat,G385gat);
nand gate_116(G462gat,G386gat,G387gat);
nand gate_117(G465gat,G388gat,G389gat);
nand gate_118(G468gat,G390gat,G391gat);
nand gate_119(G471gat,G392gat,G393gat);
nand gate_120(G474gat,G394gat,G395gat);
nand gate_121(G477gat,G396gat,G397gat);
nand gate_122(G480gat,G398gat,G399gat);
nand gate_123(G483gat,G400gat,G401gat);
nand gate_124(G486gat,G402gat,G403gat);
nand gate_125(G489gat,G404gat,G405gat);
nand gate_126(G492gat,G406gat,G407gat);
nand gate_127(G495gat,G408gat,G409gat);
nand gate_128(G498gat,G410gat,G411gat);
nand gate_129(G501gat,G412gat,G413gat);
nand gate_130(G504gat,G414gat,G415gat);
nand gate_131(G507gat,G416gat,G417gat);
nand gate_132(G510gat,G418gat,G419gat);
nand gate_133(G513gat,G420gat,G421gat);
nand gate_134(G516gat,G422gat,G423gat);
nand gate_135(G519gat,G424gat,G425gat);
nand gate_136(G522gat,G426gat,G429gat);
nand gate_137(G525gat,G432gat,G435gat);
nand gate_138(G528gat,G438gat,G441gat);
nand gate_139(G531gat,G444gat,G447gat);
nand gate_140(G534gat,G450gat,G453gat);
nand gate_141(G537gat,G456gat,G459gat);
nand gate_142(G540gat,G462gat,G465gat);
nand gate_143(G543gat,G468gat,G471gat);
nand gate_144(G546gat,G474gat,G477gat);
nand gate_145(G549gat,G480gat,G483gat);
nand gate_146(G552gat,G486gat,G489gat);
nand gate_147(G555gat,G492gat,G495gat);
nand gate_148(G558gat,G498gat,G501gat);
nand gate_149(G561gat,G504gat,G507gat);
nand gate_150(G564gat,G510gat,G513gat);
nand gate_151(G567gat,G516gat,G519gat);
nand gate_152(G570gat,G426gat,G522gat);
nand gate_153(G571gat,G429gat,G522gat);
nand gate_154(G572gat,G432gat,G525gat);
nand gate_155(G573gat,G435gat,G525gat);
nand gate_156(G574gat,G438gat,G528gat);
nand gate_157(G575gat,G441gat,G528gat);
nand gate_158(G576gat,G444gat,G531gat);
nand gate_159(G577gat,G447gat,G531gat);
nand gate_160(G578gat,G450gat,G534gat);
nand gate_161(G579gat,G453gat,G534gat);
nand gate_162(G580gat,G456gat,G537gat);
nand gate_163(G581gat,G459gat,G537gat);
nand gate_164(G582gat,G462gat,G540gat);
nand gate_165(G583gat,G465gat,G540gat);
nand gate_166(G584gat,G468gat,G543gat);
nand gate_167(G585gat,G471gat,G543gat);
nand gate_168(G586gat,G474gat,G546gat);
nand gate_169(G587gat,G477gat,G546gat);
nand gate_170(G588gat,G480gat,G549gat);
nand gate_171(G589gat,G483gat,G549gat);
nand gate_172(G590gat,G486gat,G552gat);
nand gate_173(G591gat,G489gat,G552gat);
nand gate_174(G592gat,G492gat,G555gat);
nand gate_175(G593gat,G495gat,G555gat);
nand gate_176(G594gat,G498gat,G558gat);
nand gate_177(G595gat,G501gat,G558gat);
nand gate_178(G596gat,G504gat,G561gat);
nand gate_179(G597gat,G507gat,G561gat);
nand gate_180(G598gat,G510gat,G564gat);
nand gate_181(G599gat,G513gat,G564gat);
nand gate_182(G600gat,G516gat,G567gat);
nand gate_183(G601gat,G519gat,G567gat);
nand gate_184(G602gat,G570gat,G571gat);
nand gate_185(G607gat,G572gat,G573gat);
nand gate_186(G612gat,G574gat,G575gat);
nand gate_187(G617gat,G576gat,G577gat);
nand gate_188(G622gat,G578gat,G579gat);
nand gate_189(G627gat,G580gat,G581gat);
nand gate_190(G632gat,G582gat,G583gat);
nand gate_191(G637gat,G584gat,G585gat);
nand gate_192(G642gat,G586gat,G587gat);
nand gate_193(G645gat,G588gat,G589gat);
nand gate_194(G648gat,G590gat,G591gat);
nand gate_195(G651gat,G592gat,G593gat);
nand gate_196(G654gat,G594gat,G595gat);
nand gate_197(G657gat,G596gat,G597gat);
nand gate_198(G660gat,G598gat,G599gat);
nand gate_199(G663gat,G600gat,G601gat);
nand gate_200(G666gat,G602gat,G607gat);
nand gate_201(G669gat,G612gat,G617gat);
nand gate_202(G672gat,G602gat,G612gat);
nand gate_203(G675gat,G607gat,G617gat);
nand gate_204(G678gat,G622gat,G627gat);
nand gate_205(G681gat,G632gat,G637gat);
nand gate_206(G684gat,G622gat,G632gat);
nand gate_207(G687gat,G627gat,G637gat);
nand gate_208(G690gat,G602gat,G666gat);
nand gate_209(G691gat,G607gat,G666gat);
nand gate_210(G692gat,G612gat,G669gat);
nand gate_211(G693gat,G617gat,G669gat);
nand gate_212(G694gat,G602gat,G672gat);
nand gate_213(G695gat,G612gat,G672gat);
nand gate_214(G696gat,G607gat,G675gat);
nand gate_215(G697gat,G617gat,G675gat);
nand gate_216(G698gat,G622gat,G678gat);
nand gate_217(G699gat,G627gat,G678gat);
nand gate_218(G700gat,G632gat,G681gat);
nand gate_219(G701gat,G637gat,G681gat);
nand gate_220(G702gat,G622gat,G684gat);
nand gate_221(G703gat,G632gat,G684gat);
nand gate_222(G704gat,G627gat,G687gat);
nand gate_223(G705gat,G637gat,G687gat);
nand gate_224(G706gat,G690gat,G691gat);
nand gate_225(G709gat,G692gat,G693gat);
nand gate_226(G712gat,G694gat,G695gat);
nand gate_227(G715gat,G696gat,G697gat);
nand gate_228(G718gat,G698gat,G699gat);
nand gate_229(G721gat,G700gat,G701gat);
nand gate_230(G724gat,G702gat,G703gat);
nand gate_231(G727gat,G704gat,G705gat);
nand gate_232(G730gat,G242gat,G718gat);
nand gate_233(G733gat,G245gat,G721gat);
nand gate_234(G736gat,G248gat,G724gat);
nand gate_235(G739gat,G251gat,G727gat);
nand gate_236(G742gat,G254gat,G706gat);
nand gate_237(G745gat,G257gat,G709gat);
nand gate_238(G748gat,G260gat,G712gat);
nand gate_239(G751gat,G263gat,G715gat);
nand gate_240(G754gat,G242gat,G730gat);
nand gate_241(G755gat,G718gat,G730gat);
nand gate_242(G756gat,G245gat,G733gat);
nand gate_243(G757gat,G721gat,G733gat);
nand gate_244(G758gat,G248gat,G736gat);
nand gate_245(G759gat,G724gat,G736gat);
nand gate_246(G760gat,G251gat,G739gat);
nand gate_247(G761gat,G727gat,G739gat);
nand gate_248(G762gat,G254gat,G742gat);
nand gate_249(G763gat,G706gat,G742gat);
nand gate_250(G764gat,G257gat,G745gat);
nand gate_251(G765gat,G709gat,G745gat);
nand gate_252(G766gat,G260gat,G748gat);
nand gate_253(G767gat,G712gat,G748gat);
nand gate_254(G768gat,G263gat,G751gat);
nand gate_255(G769gat,G715gat,G751gat);
nand gate_256(G770gat,G754gat,G755gat);
nand gate_257(G773gat,G756gat,G757gat);
nand gate_258(G776gat,G758gat,G759gat);
nand gate_259(G779gat,G760gat,G761gat);
nand gate_260(G782gat,G762gat,G763gat);
nand gate_261(G785gat,G764gat,G765gat);
nand gate_262(G788gat,G766gat,G767gat);
nand gate_263(G791gat,G768gat,G769gat);
nand gate_264(G794gat,G642gat,G770gat);
nand gate_265(G797gat,G645gat,G773gat);
nand gate_266(G800gat,G648gat,G776gat);
nand gate_267(G803gat,G651gat,G779gat);
nand gate_268(G806gat,G654gat,G782gat);
nand gate_269(G809gat,G657gat,G785gat);
nand gate_270(G812gat,G660gat,G788gat);
nand gate_271(G815gat,G663gat,G791gat);
nand gate_272(G818gat,G642gat,G794gat);
nand gate_273(G819gat,G770gat,G794gat);
nand gate_274(G820gat,G645gat,G797gat);
nand gate_275(G821gat,G773gat,G797gat);
nand gate_276(G822gat,G648gat,G800gat);
nand gate_277(G823gat,G776gat,G800gat);
nand gate_278(G824gat,G651gat,G803gat);
nand gate_279(G825gat,G779gat,G803gat);
nand gate_280(G826gat,G654gat,G806gat);
nand gate_281(G827gat,G782gat,G806gat);
nand gate_282(G828gat,G657gat,G809gat);
nand gate_283(G829gat,G785gat,G809gat);
nand gate_284(G830gat,G660gat,G812gat);
nand gate_285(G831gat,G788gat,G812gat);
nand gate_286(G832gat,G663gat,G815gat);
nand gate_287(G833gat,G791gat,G815gat);
nand gate_288(G834gat,G818gat,G819gat);
nand gate_289(G847gat,G820gat,G821gat);
nand gate_290(G860gat,G822gat,G823gat);
nand gate_291(G873gat,G824gat,G825gat);
nand gate_292(G886gat,G828gat,G829gat);
nand gate_293(G899gat,G832gat,G833gat);
nand gate_294(G912gat,G830gat,G831gat);
nand gate_295(G925gat,G826gat,G827gat);
not gate_296(G938gat,G834gat);
not gate_297(G939gat,G847gat);
not gate_298(G940gat,G860gat);
not gate_299(G941gat,G834gat);
not gate_300(G942gat,G847gat);
not gate_301(G943gat,G873gat);
not gate_302(G944gat,G834gat);
not gate_303(G945gat,G860gat);
not gate_304(G946gat,G873gat);
not gate_305(G947gat,G847gat);
not gate_306(G948gat,G860gat);
not gate_307(G949gat,G873gat);
not gate_308(G950gat,G886gat);
not gate_309(G951gat,G899gat);
not gate_310(G952gat,G886gat);
not gate_311(G953gat,G912gat);
not gate_312(G954gat,G925gat);
not gate_313(G955gat,G899gat);
not gate_314(G956gat,G925gat);
not gate_315(G957gat,G912gat);
not gate_316(G958gat,G925gat);
not gate_317(G959gat,G886gat);
not gate_318(G960gat,G912gat);
not gate_319(G961gat,G925gat);
not gate_320(G962gat,G886gat);
not gate_321(G963gat,G899gat);
not gate_322(G964gat,G925gat);
not gate_323(G965gat,G912gat);
not gate_324(G966gat,G899gat);
not gate_325(G967gat,G886gat);
not gate_326(G968gat,G912gat);
not gate_327(G969gat,G899gat);
not gate_328(G970gat,G847gat);
not gate_329(G971gat,G873gat);
not gate_330(G972gat,G847gat);
not gate_331(G973gat,G860gat);
not gate_332(G974gat,G834gat);
not gate_333(G975gat,G873gat);
not gate_334(G976gat,G834gat);
not gate_335(G977gat,G860gat);
and gate_336(G978gat,G938gat,G939gat,G940gat,G873gat);
and gate_337(G979gat,G941gat,G942gat,G860gat,G943gat);
and gate_338(G980gat,G944gat,G847gat,G945gat,G946gat);
and gate_339(G981gat,G834gat,G947gat,G948gat,G949gat);
and gate_340(G982gat,G958gat,G959gat,G960gat,G899gat);
and gate_341(G983gat,G961gat,G962gat,G912gat,G963gat);
and gate_342(G984gat,G964gat,G886gat,G965gat,G966gat);
and gate_343(G985gat,G925gat,G967gat,G968gat,G969gat);
or gate_344(G986gat,G978gat,G979gat,G980gat,G981gat);
or gate_345(G991gat,G982gat,G983gat,G984gat,G985gat);
and gate_346(G996gat,G925gat,G950gat,G912gat,G951gat,G986gat);
and gate_347(G1001gat,G925gat,G952gat,G953gat,G899gat,G986gat);
and gate_348(G1006gat,G954gat,G886gat,G912gat,G955gat,G986gat);
and gate_349(G1011gat,G956gat,G886gat,G957gat,G899gat,G986gat);
and gate_350(G1016gat,G834gat,G970gat,G860gat,G971gat,G991gat);
and gate_351(G1021gat,G834gat,G972gat,G973gat,G873gat,G991gat);
and gate_352(G1026gat,G974gat,G847gat,G860gat,G975gat,G991gat);
and gate_353(G1031gat,G976gat,G847gat,G977gat,G873gat,G991gat);
and gate_354(G1036gat,G834gat,G996gat);
and gate_355(G1039gat,G847gat,G996gat);
and gate_356(G1042gat,G860gat,G996gat);
and gate_357(G1045gat,G873gat,G996gat);
and gate_358(G1048gat,G834gat,G1001gat);
and gate_359(G1051gat,G847gat,G1001gat);
and gate_360(G1054gat,G860gat,G1001gat);
and gate_361(G1057gat,G873gat,G1001gat);
and gate_362(G1060gat,G834gat,G1006gat);
and gate_363(G1063gat,G847gat,G1006gat);
and gate_364(G1066gat,G860gat,G1006gat);
and gate_365(G1069gat,G873gat,G1006gat);
and gate_366(G1072gat,G834gat,G1011gat);
and gate_367(G1075gat,G847gat,G1011gat);
and gate_368(G1078gat,G860gat,G1011gat);
and gate_369(G1081gat,G873gat,G1011gat);
and gate_370(G1084gat,G925gat,G1016gat);
and gate_371(G1087gat,G886gat,G1016gat);
and gate_372(G1090gat,G912gat,G1016gat);
and gate_373(G1093gat,G899gat,G1016gat);
and gate_374(G1096gat,G925gat,G1021gat);
and gate_375(G1099gat,G886gat,G1021gat);
and gate_376(G1102gat,G912gat,G1021gat);
and gate_377(G1105gat,G899gat,G1021gat);
and gate_378(G1108gat,G925gat,G1026gat);
and gate_379(G1111gat,G886gat,G1026gat);
and gate_380(G1114gat,G912gat,G1026gat);
and gate_381(G1117gat,G899gat,G1026gat);
and gate_382(G1120gat,G925gat,G1031gat);
and gate_383(G1123gat,G886gat,G1031gat);
and gate_384(G1126gat,G912gat,G1031gat);
and gate_385(G1129gat,G899gat,G1031gat);
nand gate_386(G1132gat,G1gat,G1036gat);
nand gate_387(G1135gat,G8gat,G1039gat);
nand gate_388(G1138gat,G15gat,G1042gat);
nand gate_389(G1141gat,G22gat,G1045gat);
nand gate_390(G1144gat,G29gat,G1048gat);
nand gate_391(G1147gat,G36gat,G1051gat);
nand gate_392(G1150gat,G43gat,G1054gat);
nand gate_393(G1153gat,G50gat,G1057gat);
nand gate_394(G1156gat,G57gat,G1060gat);
nand gate_395(G1159gat,G64gat,G1063gat);
nand gate_396(G1162gat,G71gat,G1066gat);
nand gate_397(G1165gat,G78gat,G1069gat);
nand gate_398(G1168gat,G85gat,G1072gat);
nand gate_399(G1171gat,G92gat,G1075gat);
nand gate_400(G1174gat,G99gat,G1078gat);
nand gate_401(G1177gat,G106gat,G1081gat);
nand gate_402(G1180gat,G113gat,G1084gat);
nand gate_403(G1183gat,G120gat,G1087gat);
nand gate_404(G1186gat,G127gat,G1090gat);
nand gate_405(G1189gat,G134gat,G1093gat);
nand gate_406(G1192gat,G141gat,G1096gat);
nand gate_407(G1195gat,G148gat,G1099gat);
nand gate_408(G1198gat,G155gat,G1102gat);
nand gate_409(G1201gat,G162gat,G1105gat);
nand gate_410(G1204gat,G169gat,G1108gat);
nand gate_411(G1207gat,G176gat,G1111gat);
nand gate_412(G1210gat,G183gat,G1114gat);
nand gate_413(G1213gat,G190gat,G1117gat);
nand gate_414(G1216gat,G197gat,G1120gat);
nand gate_415(G1219gat,G204gat,G1123gat);
nand gate_416(G1222gat,G211gat,G1126gat);
nand gate_417(G1225gat,G218gat,G1129gat);
nand gate_418(G1228gat,G1gat,G1132gat);
nand gate_419(G1229gat,G1036gat,G1132gat);
nand gate_420(G1230gat,G8gat,G1135gat);
nand gate_421(G1231gat,G1039gat,G1135gat);
nand gate_422(G1232gat,G15gat,G1138gat);
nand gate_423(G1233gat,G1042gat,G1138gat);
nand gate_424(G1234gat,G22gat,G1141gat);
nand gate_425(G1235gat,G1045gat,G1141gat);
nand gate_426(G1236gat,G29gat,G1144gat);
nand gate_427(G1237gat,G1048gat,G1144gat);
nand gate_428(G1238gat,G36gat,G1147gat);
nand gate_429(G1239gat,G1051gat,G1147gat);
nand gate_430(G1240gat,G43gat,G1150gat);
nand gate_431(G1241gat,G1054gat,G1150gat);
nand gate_432(G1242gat,G50gat,G1153gat);
nand gate_433(G1243gat,G1057gat,G1153gat);
nand gate_434(G1244gat,G57gat,G1156gat);
nand gate_435(G1245gat,G1060gat,G1156gat);
nand gate_436(G1246gat,G64gat,G1159gat);
nand gate_437(G1247gat,G1063gat,G1159gat);
nand gate_438(G1248gat,G71gat,G1162gat);
nand gate_439(G1249gat,G1066gat,G1162gat);
nand gate_440(G1250gat,G78gat,G1165gat);
nand gate_441(G1251gat,G1069gat,G1165gat);
nand gate_442(G1252gat,G85gat,G1168gat);
nand gate_443(G1253gat,G1072gat,G1168gat);
nand gate_444(G1254gat,G92gat,G1171gat);
nand gate_445(G1255gat,G1075gat,G1171gat);
nand gate_446(G1256gat,G99gat,G1174gat);
nand gate_447(G1257gat,G1078gat,G1174gat);
nand gate_448(G1258gat,G106gat,G1177gat);
nand gate_449(G1259gat,G1081gat,G1177gat);
nand gate_450(G1260gat,G113gat,G1180gat);
nand gate_451(G1261gat,G1084gat,G1180gat);
nand gate_452(G1262gat,G120gat,G1183gat);
nand gate_453(G1263gat,G1087gat,G1183gat);
nand gate_454(G1264gat,G127gat,G1186gat);
nand gate_455(G1265gat,G1090gat,G1186gat);
nand gate_456(G1266gat,G134gat,G1189gat);
nand gate_457(G1267gat,G1093gat,G1189gat);
nand gate_458(G1268gat,G141gat,G1192gat);
nand gate_459(G1269gat,G1096gat,G1192gat);
nand gate_460(G1270gat,G148gat,G1195gat);
nand gate_461(G1271gat,G1099gat,G1195gat);
nand gate_462(G1272gat,G155gat,G1198gat);
nand gate_463(G1273gat,G1102gat,G1198gat);
nand gate_464(G1274gat,G162gat,G1201gat);
nand gate_465(G1275gat,G1105gat,G1201gat);
nand gate_466(G1276gat,G169gat,G1204gat);
nand gate_467(G1277gat,G1108gat,G1204gat);
nand gate_468(G1278gat,G176gat,G1207gat);
nand gate_469(G1279gat,G1111gat,G1207gat);
nand gate_470(G1280gat,G183gat,G1210gat);
nand gate_471(G1281gat,G1114gat,G1210gat);
nand gate_472(G1282gat,G190gat,G1213gat);
nand gate_473(G1283gat,G1117gat,G1213gat);
nand gate_474(G1284gat,G197gat,G1216gat);
nand gate_475(G1285gat,G1120gat,G1216gat);
nand gate_476(G1286gat,G204gat,G1219gat);
nand gate_477(G1287gat,G1123gat,G1219gat);
nand gate_478(G1288gat,G211gat,G1222gat);
nand gate_479(G1289gat,G1126gat,G1222gat);
nand gate_480(G1290gat,G218gat,G1225gat);
nand gate_481(G1291gat,G1129gat,G1225gat);
nand gate_482(G1292gat,G1228gat,G1229gat);
nand gate_483(G1293gat,G1230gat,G1231gat);
nand gate_484(G1294gat,G1232gat,G1233gat);
nand gate_485(G1295gat,G1234gat,G1235gat);
nand gate_486(G1296gat,G1236gat,G1237gat);
nand gate_487(G1297gat,G1238gat,G1239gat);
nand gate_488(G1298gat,G1240gat,G1241gat);
nand gate_489(G1299gat,G1242gat,G1243gat);
nand gate_490(G1300gat,G1244gat,G1245gat);
nand gate_491(G1301gat,G1246gat,G1247gat);
nand gate_492(G1302gat,G1248gat,G1249gat);
nand gate_493(G1303gat,G1250gat,G1251gat);
nand gate_494(G1304gat,G1252gat,G1253gat);
nand gate_495(G1305gat,G1254gat,G1255gat);
nand gate_496(G1306gat,G1256gat,G1257gat);
nand gate_497(G1307gat,G1258gat,G1259gat);
nand gate_498(G1308gat,G1260gat,G1261gat);
nand gate_499(G1309gat,G1262gat,G1263gat);
nand gate_500(G1310gat,G1264gat,G1265gat);
nand gate_501(G1311gat,G1266gat,G1267gat);
nand gate_502(G1312gat,G1268gat,G1269gat);
nand gate_503(G1313gat,G1270gat,G1271gat);
nand gate_504(G1314gat,G1272gat,G1273gat);
nand gate_505(G1315gat,G1274gat,G1275gat);
nand gate_506(G1316gat,G1276gat,G1277gat);
nand gate_507(G1317gat,G1278gat,G1279gat);
nand gate_508(G1318gat,G1280gat,G1281gat);
nand gate_509(G1319gat,G1282gat,G1283gat);
nand gate_510(G1320gat,G1284gat,G1285gat);
nand gate_511(G1321gat,G1286gat,G1287gat);
nand gate_512(G1322gat,G1288gat,G1289gat);
nand gate_513(G1323gat,G1290gat,G1291gat);
buf gate_514(G1324gat,G1292gat);
buf gate_515(G1325gat,G1293gat);
buf gate_516(G1326gat,G1294gat);
buf gate_517(G1327gat,G1295gat);
buf gate_518(G1328gat,G1296gat);
buf gate_519(G1329gat,G1297gat);
buf gate_520(G1330gat,G1298gat);
buf gate_521(G1331gat,G1299gat);
buf gate_522(G1332gat,G1300gat);
buf gate_523(G1333gat,G1301gat);
buf gate_524(G1334gat,G1302gat);
buf gate_525(G1335gat,G1303gat);
buf gate_526(G1336gat,G1304gat);
buf gate_527(G1337gat,G1305gat);
buf gate_528(G1338gat,G1306gat);
buf gate_529(G1339gat,G1307gat);
buf gate_530(G1340gat,G1308gat);
buf gate_531(G1341gat,G1309gat);
buf gate_532(G1342gat,G1310gat);
buf gate_533(G1343gat,G1311gat);
buf gate_534(G1344gat,G1312gat);
buf gate_535(G1345gat,G1313gat);
buf gate_536(G1346gat,G1314gat);
buf gate_537(G1347gat,G1315gat);
buf gate_538(G1348gat,G1316gat);
buf gate_539(G1349gat,G1317gat);
buf gate_540(G1350gat,G1318gat);
buf gate_541(G1351gat,G1319gat);
buf gate_542(G1352gat,G1320gat);
buf gate_543(G1353gat,G1321gat);
buf gate_544(G1354gat,G1322gat);
buf gate_545(G1355gat,G1323gat);
endmodule
