// Verilog File 
module k2 (vdd,pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,
pi08,pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,
pi18,pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,
pi28,pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,
pi38,pi39,pi40,pi41,pi42,pi43,pi44,po00,po01,po02,
po03,po04,po05,po06,po07,po08,po09,po10,po11,po12,
po13,po14,po15,po16,po17,po18,po19,po20,po21,po22,
po23,po24,po25,po26,po27,po28,po29,po30,po31,po32,
po33,po34,po35,po36,po37,po38,po39,po40,po41,po42,
po43,po44);

input vdd,pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,
pi08,pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,
pi18,pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,
pi28,pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,
pi38,pi39,pi40,pi41,pi42,pi43,pi44;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18,
po19,po20,po21,po22,po23,po24,po25,po26,po27,po28,
po29,po30,po31,po32,po33,po34,po35,po36,po37,po38,
po39,po40,po41,po42,po43,po44;

wire n90,n92,n93,n94,n95,n96,n97,n98,n99,
n100,n101,n102,n103,n104,n105,n106,n107,n108,n109,
n110,n111,n112,n113,n114,n115,n116,n117,n118,n119,
n120,n121,n122,n123,n124,n125,n126,n127,n128,n129,
n130,n131,n132,n133,n134,n135,n136,n137,n138,n139,
n140,n141,n142,n143,n144,n145,n146,n147,n148,n149,
n150,n151,n152,n153,n154,n155,n156,n157,n158,n159,
n160,n161,n162,n163,n164,n165,n166,n167,n168,n170,
n171,n172,n173,n174,n175,n176,n177,n178,n180,n182,
n184,n185,n186,n187,n188,n189,n190,n191,n192,n193,
n194,n195,n196,n197,n198,n199,n200,n201,n202,n203,
n204,n205,n206,n207,n209,n210,n211,n212,n213,n214,
n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,
n225,n226,n227,n228,n229,n230,n231,n232,n233,n234,
n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,
n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,
n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,
n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,
n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,
n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,
n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,
n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,
n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,
n325,n326,n327,n328,n329,n330,n331,n332,n333,n334,
n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,
n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,
n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,
n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,
n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,
n385,n386,n387,n388,n389,n390,n391,n392,n393,n394,
n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,
n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,
n415,n416,n417,n418,n419,n420,n421,n422,n424,n425,
n426,n427,n428,n429,n431,n432,n433,n434,n435,n437,
n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,
n448,n450,n452,n453,n454,n455,n456,n457,n458,n459,
n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,
n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,
n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,
n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,
n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,
n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,
n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,
n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,
n540,n541,n542,n544,n545,n547,n548,n549,n550,n551,
n552,n553,n554,n555,n556,n557,n558,n559,n560,n561,
n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,
n572,n573,n574,n575,n576,n577,n578,n579,n580,n581,
n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,
n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,
n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,
n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,
n622,n623,n624,n625,n626,n627,n628,n629,n630,n631,
n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,
n642,n643,n644,n645,n646,n647,n648,n649,n650,n651,
n652,n653,n654,n655,n656,n658,n659,n660,n661,n662,
n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,
n673,n674,n675,n676,n677,n678,n679,n680,n681,n682,
n683,n684,n685,n686,n687,n688,n689,n690,n691,n692,
n693,n694,n695,n696,n697,n698,n699,n700,n701,n702,
n703,n704,n705,n706,n707,n708,n709,n710,n711,n712,
n713,n714,n715,n716,n717,n719,n720,n721,n722,n723,
n724,n725,n726,n727,n728,n729,n730,n731,n732,n733,
n734,n735,n736,n737,n738,n739,n740,n741,n742,n743,
n744,n745,n746,n747,n748,n749,n750,n751,n752,n753,
n754,n755,n756,n757,n758,n759,n760,n762,n763,n764,
n765,n766,n767,n768,n769,n770,n771,n772,n773,n774,
n775,n776,n777,n778,n779,n780,n781,n782,n783,n784,
n785,n786,n787,n788,n789,n790,n791,n792,n793,n794,
n795,n796,n797,n798,n799,n800,n801,n802,n803,n804,
n805,n806,n807,n808,n809,n810,n811,n812,n813,n814,
n815,n816,n817,n818,n819,n820,n821,n822,n823,n824,
n825,n826,n827,n828,n829,n830,n831,n832,n833,n834,
n835,n836,n837,n838,n839,n840,n841,n842,n843,n844,
n845,n846,n847,n848,n849,n850,n851,n852,n853,n854,
n855,n856,n857,n858,n859,n860,n862,n863,n864,n865,
n866,n867,n868,n869,n870,n871,n872,n873,n874,n875,
n876,n877,n878,n879,n880,n881,n882,n883,n884,n885,
n886,n887,n888,n889,n890,n891,n892,n893,n894,n895,
n897,n898,n899,n900,n901,n902,n903,n904,n905,n906,
n907,n908,n909,n910,n911,n912,n913,n914,n915,n916,
n917,n918,n919,n920,n921,n922,n923,n924,n925,n926,
n927,n928,n929,n930,n931,n932,n933,n934,n935,n936,
n937,n938,n939,n940,n941,n942,n943,n944,n945,n946,
n947,n948,n949,n950,n951,n952,n953,n954,n955,n956,
n957,n958,n959,n960,n961,n962,n963,n964,n965,n966,
n967,n968,n969,n970,n971,n972,n973,n974,n975,n976,
n977,n978,n979,n980,n981,n982,n983,n984,n985,n986,
n987,n988,n989,n990,n991,n992,n993,n994,n995,n996,
n997,n998,n999,n1000,n1001,n1002,n1003,n1004,n1005,n1006,
n1007,n1008,n1009,n1010,n1011,n1012,n1013,n1014,n1015,n1016,
n1017,n1018,n1019,n1021,n1022,n1023,n1024,n1025,n1026,n1027,
n1028,n1029,n1030,n1031,n1032,n1033,n1034,n1035,n1036,n1037,
n1038,n1039,n1040,n1041,n1042,n1043,n1044,n1045,n1046,n1047,
n1048,n1049,n1050,n1052,n1053,n1054,n1055,n1056,n1057,n1058,
n1059,n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,
n1069,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,n1079,
n1080,n1081,n1082,n1083,n1084,n1085,n1086,n1087,n1088,n1089,
n1090,n1091,n1092,n1093,n1094,n1095,n1096,n1097,n1098,n1099,
n1100,n1101,n1102,n1103,n1104,n1105,n1106,n1107,n1108,n1109,
n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,n1118,n1119,
n1120,n1121,n1123,n1124,n1125,n1126,n1127,n1128,n1129,n1130,
n1131,n1132,n1133,n1134,n1135,n1136,n1137,n1138,n1139,n1140,
n1141,n1142,n1143,n1144,n1145,n1146,n1147,n1148,n1149,n1150,
n1151,n1152,n1153,n1154,n1155,n1157,n1158,n1159,n1160,n1161,
n1162,n1163,n1164,n1165,n1166,n1167,n1168,n1169,n1170,n1171,
n1172,n1173,n1174,n1175,n1176,n1177,n1178,n1179,n1180,n1181,
n1182,n1183,n1184,n1185,n1186,n1187,n1188,n1189,n1190,n1191,
n1193,n1194,n1195,n1196,n1197,n1198,n1199,n1200,n1201,n1202,
n1203,n1204,n1205,n1206,n1207,n1208,n1209,n1210,n1211,n1212,
n1213,n1214,n1215,n1216,n1217,n1218,n1219,n1220,n1221,n1222,
n1223,n1224,n1225,n1226,n1227,n1228,n1229,n1230,n1231,n1232,
n1233,n1234,n1235,n1236,n1237,n1238,n1239,n1240,n1241,n1242,
n1243,n1244,n1245,n1246,n1247,n1248,n1249,n1250,n1251,n1252,
n1253,n1254,n1255,n1256,n1257,n1258,n1259,n1260,n1261,n1262,
n1263,n1264,n1265,n1266,n1267,n1268,n1269,n1270,n1271,n1272,
n1273,n1274,n1275,n1276,n1277,n1278,n1279,n1280,n1281,n1282,
n1283,n1284,n1285,n1286,n1287,n1288,n1289,n1290,n1291,n1292,
n1293,n1294,n1295,n1296,n1297,n1299,n1301,n1302,n1303,n1304,
n1305,n1306,n1307,n1308,n1309,n1310,n1311,n1312,n1313,n1314,
n1315,n1316,n1318,n1319,n1320,n1321,n1322,n1323,n1324,n1325,
n1326,n1327,n1328,n1329,n1330,n1331,n1332,n1333,n1334,n1335,
n1337,n1338,n1339,n1341,n1342,n1343,n1344,n1345,n1346,n1347,
n1349,n1350,n1351,n1352,n1353,n1354,n1355,n1356,n1357,n1358,
n1359,n1360,n1361,n1362,n1363,n1364,n1365,n1366,n1367,n1368,
n1369,n1370,n1371,n1372,n1373,n1374,n1375,n1376,n1377,n1378,
n1379,n1380,n1381,n1382,n1383,n1384,n1385,n1386,n1387,n1388,
n1389,n1390,n1391,n1392,n1393,n1394,n1395,n1396,n1397,n1398,
n1399,n1400,n1401,n1402,n1403,n1404,n1405,n1406,n1407,n1409,
n1410,n1411,n1412,n1413,n1414,n1415,n1416,n1417,n1418,n1419,
n1420,n1421,n1422,n1423,n1424,n1425,n1426,n1427,n1429,n1430,
n1431,n1432,n1434,n1435,n1436,n1438,n1439,n1440,n1441,n1442,
n1444,n1445,n1446,n1448,n1449,n1450,n1451,n1452,n1453,n1454,
n1455,n1456,n1457,n1458,n1459,n1460,n1461,n1462,n1463,n1464,
n1465,n1466,n1467,n1468,n1469,n1470,n1471,n1472,n1473,n1474,
n1475,n1476,n1477,n1478,n1479,n1480,n1481,n1482,n1483,n1484,
n1485,n1486,n1487,n1488,n1489,n1490,n1491,n1492,n1493,n1494,
n1495,n1497,n1498,n1499,n1500,n1501,n1502,n1503,n1504,n1505,
n1506,n1507,n1508,n1509,n1510,n1511,n1512,n1513,n1514,n1515,
n1516,n1517,n1518,n1519,n1520,n1521,n1522,n1523,n1524,n1525,
n1526,n1527,n1528,n1529,n1530,n1531,n1532,n1533,n1534,n1535,
n1536,n1537,n1538,n1539,n1540,n1541,n1542,n1543,n1544,n1545,
n1546,n1547,n1548,n1549,n1550,n1551,n1552,n1553,n1554,n1555,
n1556,n1557,n1558,n1559,n1560,n1561,n1562,n1563,n1564,n1566,
n1567,n1568,n1569,n1570,n1571,n1572,n1573,n1574,n1575,n1576,
n1577,n1578,n1579,n1580,n1581,n1582,n1583,n1584,n1585,n1586,
n1587,n1588,n1589,n1590,n1591,n1592,n1593,n1594,n1595,n1596,
n1597,n1598,n1599,n1600,n1601,n1602,n1603,n1604,n1605,n1606,
n1607,n1608,n1609,n1610,n1611,n1612,n1613,n1614,n1615,n1616,
n1617,n1618,n1619,n1620,n1621,n1622,n1623,n1624,n1625,n1626,
n1627,n1628,n1629,n1630,n1631,n1632,n1633,n1634,n1635,n1636,
n1637,n1638,n1639,n1640,n1641,n1642,n1643,n1644,n1645,n1646,
n1647,n1648,n1649,n1650,n1651,n1652,n1653,n1655,n1656,n1657,
n1658,n1659,n1660,n1661,n1662,n1663,n1664,n1665,n1666,n1667,
n1668,n1669,n1670,n1671,n1672,n1673,n1674,n1675,n1676,n1677,
n1678,n1679,n1680,n1681,n1682,n1683,n1684,n1685,n1686,n1687,
n1688,n1689,n1690,n1691,n1692,n1693,n1694,n1695,n1696,n1697,
n1698,n1699,n1700,n1701,n1702,n1703,n1704,n1705,n1706,n1707,
n1708,n1709,n1710,n1711,n1712,n1713,n1714,n1715,n1716,n1717,
n1718,n1719,n1720,n1721,n1722,n1723,n1724,n1725,n1726,n1727,
n1728,n1729,n1730,n1731,n1732,n1733,n1734,n1735,n1736,n1737,
n1738,n1739,n1740,n1741,n1742,n1743,n1744,n1745,n1746,n1747,
n1748,n1749,n1750,n1751,n1752,n1753,n1754,n1755,n1756,n1757,
n1758,n1759,n1760,n1762,n1763,n1764,n1765,n1766,n1767,n1768,
n1769,n1770,n1771,n1772,n1773,n1774,n1775,n1776,n1777,n1778,
n1779,n1780,n1781,n1782,n1783,n1784,n1785,n1786,n1787,n1788,
n1789,n1790,n1791,n1792,n1793,n1794,n1795,n1796,n1797,n1798,
n1799,n1800,n1801,n1802,n1803,n1804,n1805,n1806,n1807,n1808,
n1809,n1810,n1811,n1812,n1813,n1814,n1815,n1816,n1817,n1818,
n1819,n1820,n1821,n1822,n1823,n1824,n1825,n1826,n1827,n1828,
n1829,n1830,n1831,n1832,n1833,n1834,n1835,n1836,n1837,n1838,
n1839,n1840,n1841,n1842,n1843,n1844,n1845,n1846,n1847,n1848,
n1849,n1850,n1851,n1852,n1853,n1854,n1855,n1856,n1857,n1858,
n1859,n1860,n1861,n1862,n1863,n1864,n1865,n1866,n1867,n1868,
n1869,n1870,n1871,n1872,n1873,n1874,n1875,n1876,n1877,n1878,
n1879,n1880,n1881,n1882,n1883,n1884,n1886,n1887,n1888,n1889,
n1890,n1891,n1892,n1893,n1894,n1895,n1897,n1898,n1899,n1900,
n1901;
buf gate_0(n90,vdd);
not gate_1(po02,n90);
not gate_2(n92,pi00);
not gate_3(n93,pi01);
not gate_4(n94,pi02);
not gate_5(n95,pi03);
not gate_6(n96,pi04);
not gate_7(n97,pi05);
not gate_8(n98,pi06);
not gate_9(n99,pi07);
not gate_10(n100,pi08);
not gate_11(n101,pi09);
not gate_12(n102,pi10);
not gate_13(n103,pi11);
not gate_14(n104,pi12);
not gate_15(n105,pi13);
not gate_16(n106,pi14);
not gate_17(n107,pi15);
not gate_18(n108,pi16);
not gate_19(n109,pi17);
not gate_20(n110,pi18);
not gate_21(n111,pi19);
not gate_22(n112,pi20);
not gate_23(n113,pi21);
not gate_24(n114,pi22);
not gate_25(n115,pi23);
not gate_26(n116,pi25);
not gate_27(n117,pi26);
not gate_28(n118,pi27);
not gate_29(n119,pi28);
not gate_30(n120,pi29);
not gate_31(n121,pi30);
not gate_32(n122,pi31);
not gate_33(n123,pi32);
not gate_34(n124,pi33);
not gate_35(n125,pi34);
not gate_36(n126,pi35);
not gate_37(n127,pi36);
not gate_38(n128,pi38);
not gate_39(n129,pi39);
not gate_40(n130,pi40);
not gate_41(n131,pi41);
not gate_42(n132,pi42);
not gate_43(n133,pi43);
not gate_44(n134,pi44);
and gate_45(n135,n110,pi19);
and gate_46(n136,pi21,n135);
and gate_47(n137,pi24,n136);
and gate_48(n138,n119,n137);
and gate_49(n139,n120,pi30);
and gate_50(n140,n138,n139);
not gate_51(n141,n140);
and gate_52(n142,pi26,n119);
not gate_53(n143,n142);
and gate_54(n144,n136,n142);
and gate_55(n145,n139,n144);
not gate_56(n146,n145);
and gate_57(n147,n141,n146);
and gate_58(n148,pi10,n136);
and gate_59(n149,pi25,n148);
and gate_60(n150,n119,n149);
and gate_61(n151,n139,n150);
not gate_62(n152,n151);
and gate_63(n153,n147,n152);
and gate_64(n154,n111,pi20);
and gate_65(n155,n110,n154);
and gate_66(n156,n92,n155);
and gate_67(n157,pi21,n156);
and gate_68(n158,pi24,n157);
and gate_69(n159,n139,n158);
not gate_70(n160,n159);
and gate_71(n161,pi19,pi20);
and gate_72(n162,pi18,n161);
and gate_73(n163,n92,n162);
and gate_74(n164,pi21,n163);
and gate_75(n165,pi24,n164);
and gate_76(n166,n139,n165);
not gate_77(n167,n166);
and gate_78(n168,n160,n167);
not gate_79(po01,n168);
and gate_80(n170,pi18,n111);
and gate_81(n171,n112,n170);
and gate_82(n172,pi21,n171);
and gate_83(n173,n119,n172);
and gate_84(n174,n92,n173);
and gate_85(n175,n139,n174);
not gate_86(n176,n175);
and gate_87(n177,n168,n176);
and gate_88(n178,n153,n177);
not gate_89(po00,n178);
and gate_90(n180,n146,n152);
not gate_91(po03,n180);
and gate_92(n182,n147,n167);
not gate_93(po04,n182);
and gate_94(n184,pi00,n110);
and gate_95(n185,n154,n184);
and gate_96(n186,pi21,n185);
and gate_97(n187,pi24,n186);
and gate_98(n188,n139,n187);
not gate_99(n189,n188);
and gate_100(n190,pi19,n184);
and gate_101(n191,pi21,n190);
and gate_102(n192,pi28,n139);
not gate_103(n193,n192);
and gate_104(n194,n191,n192);
not gate_105(n195,n194);
and gate_106(n196,n189,n195);
and gate_107(n197,pi00,n173);
and gate_108(n198,n139,n197);
not gate_109(n199,n198);
and gate_110(n200,pi00,pi18);
and gate_111(n201,pi19,n200);
and gate_112(n202,pi20,n201);
and gate_113(n203,pi21,n139);
and gate_114(n204,n202,n203);
not gate_115(n205,n204);
and gate_116(n206,n199,n205);
and gate_117(n207,n196,n206);
not gate_118(po05,n207);
and gate_119(n209,pi03,pi27);
and gate_120(n210,n113,n202);
and gate_121(n211,n209,n210);
and gate_122(n212,n120,n211);
and gate_123(n213,n121,n212);
not gate_124(n214,n213);
and gate_125(n215,pi00,n97);
and gate_126(n216,pi18,pi19);
and gate_127(n217,pi20,n216);
and gate_128(n218,n113,n217);
and gate_129(n219,n118,n218);
and gate_130(n220,n119,n219);
and gate_131(n221,pi29,n220);
and gate_132(n222,n215,n221);
and gate_133(n223,pi30,n222);
not gate_134(n224,n223);
and gate_135(n225,n92,n96);
and gate_136(n226,pi28,n219);
and gate_137(n227,pi29,n226);
and gate_138(n228,n225,n227);
and gate_139(n229,n121,n228);
not gate_140(n230,n229);
and gate_141(n231,n224,n230);
and gate_142(n232,n214,n231);
and gate_143(n233,pi00,pi11);
and gate_144(n234,pi18,n233);
and gate_145(n235,pi19,n112);
and gate_146(n236,n234,n235);
and gate_147(n237,n113,n236);
and gate_148(n238,pi26,n237);
and gate_149(n239,n192,n238);
not gate_150(n240,n239);
and gate_151(n241,pi00,n103);
and gate_152(n242,pi18,n241);
and gate_153(n243,n235,n242);
and gate_154(n244,n113,n243);
and gate_155(n245,pi26,n244);
and gate_156(n246,n192,n245);
not gate_157(n247,n246);
and gate_158(n248,n240,n247);
and gate_159(n249,pi00,pi10);
and gate_160(n250,n103,n249);
and gate_161(n251,n112,n216);
and gate_162(n252,n113,n251);
and gate_163(n253,pi25,n252);
and gate_164(n254,pi29,n253);
and gate_165(n255,n250,n254);
and gate_166(n256,n121,n255);
not gate_167(n257,n256);
and gate_168(n258,pi29,n121);
and gate_169(n259,n112,n201);
and gate_170(n260,n113,n259);
and gate_171(n261,n142,n260);
and gate_172(n262,n258,n261);
not gate_173(n263,n262);
and gate_174(n264,n257,n263);
and gate_175(n265,n248,n264);
and gate_176(n266,n232,n265);
and gate_177(n267,pi22,n260);
and gate_178(n268,n258,n267);
not gate_179(n269,n268);
and gate_180(n270,pi11,n249);
and gate_181(n271,pi18,n270);
and gate_182(n272,n235,n271);
and gate_183(n273,n113,n272);
and gate_184(n274,pi25,n273);
and gate_185(n275,n258,n274);
not gate_186(n276,n275);
and gate_187(n277,n269,n276);
and gate_188(n278,n154,n242);
and gate_189(n279,n113,n278);
and gate_190(n280,pi26,n279);
and gate_191(n281,n192,n280);
not gate_192(n282,n281);
and gate_193(n283,n154,n234);
and gate_194(n284,n113,n283);
and gate_195(n285,pi26,n284);
and gate_196(n286,n192,n285);
not gate_197(n287,n286);
and gate_198(n288,n282,n287);
and gate_199(n289,n277,n288);
and gate_200(n290,pi18,n154);
and gate_201(n291,n109,n290);
and gate_202(n292,n113,n291);
and gate_203(n293,pi26,n292);
and gate_204(n294,n119,n293);
and gate_205(n295,pi29,n294);
and gate_206(n296,pi00,n295);
and gate_207(n297,n121,n296);
not gate_208(n298,n297);
and gate_209(n299,pi20,n170);
and gate_210(n300,n113,n299);
and gate_211(n301,pi26,n300);
and gate_212(n302,pi17,n301);
and gate_213(n303,n119,n302);
and gate_214(n304,pi29,n303);
and gate_215(n305,n121,n304);
not gate_216(n306,n305);
and gate_217(n307,pi00,n305);
not gate_218(n308,n307);
and gate_219(n309,n298,n308);
and gate_220(n310,n110,n215);
and gate_221(n311,n161,n310);
and gate_222(n312,n113,n311);
and gate_223(n313,pi22,n312);
and gate_224(n314,n119,n258);
not gate_225(n315,n314);
and gate_226(n316,n313,n314);
not gate_227(n317,n316);
and gate_228(n318,pi20,pi22);
and gate_229(n319,n113,n190);
and gate_230(n320,n318,n319);
and gate_231(n321,pi28,n320);
and gate_232(n322,n258,n321);
not gate_233(n323,n322);
and gate_234(n324,n317,n323);
and gate_235(n325,n309,n324);
and gate_236(n326,n289,n325);
and gate_237(n327,n266,n326);
and gate_238(n328,pi02,n95);
and gate_239(n329,n184,n328);
and gate_240(n330,n111,n329);
and gate_241(n331,n112,n330);
and gate_242(n332,n113,n331);
and gate_243(n333,n192,n332);
not gate_244(n334,n333);
and gate_245(n335,n113,n185);
and gate_246(n336,pi23,n119);
and gate_247(n337,n335,n336);
and gate_248(n338,n258,n337);
not gate_249(n339,n338);
and gate_250(n340,n334,n339);
and gate_251(n341,n94,n95);
and gate_252(n342,n110,n341);
and gate_253(n343,n111,n342);
and gate_254(n344,pi00,n343);
and gate_255(n345,pi20,n344);
and gate_256(n346,n113,n345);
and gate_257(n347,n192,n346);
not gate_258(n348,n347);
and gate_259(n349,n340,n348);
and gate_260(n350,pi21,n299);
and gate_261(n351,n97,n107);
and gate_262(n352,n241,n351);
and gate_263(n353,n350,n352);
and gate_264(n354,n142,n353);
and gate_265(n355,n139,n354);
not gate_266(n356,n355);
and gate_267(n357,pi21,n119);
and gate_268(n358,n139,n357);
not gate_269(n359,n358);
and gate_270(n360,n283,n351);
and gate_271(n361,pi26,n360);
and gate_272(n362,n358,n361);
not gate_273(n363,n362);
and gate_274(n364,n356,n363);
and gate_275(n365,n271,n351);
and gate_276(n366,n154,n365);
and gate_277(n367,pi25,n366);
and gate_278(n368,n358,n367);
not gate_279(n369,n368);
and gate_280(n370,n95,n310);
and gate_281(n371,n111,n370);
and gate_282(n372,n112,n371);
and gate_283(n373,n113,n372);
and gate_284(n374,n314,n373);
not gate_285(n375,n374);
and gate_286(n376,n369,n375);
and gate_287(n377,n364,n376);
and gate_288(n378,n349,n377);
and gate_289(n379,pi22,n186);
and gate_290(n380,n139,n379);
not gate_291(n381,n380);
and gate_292(n382,n155,n250);
and gate_293(n383,pi21,n382);
and gate_294(n384,pi25,n383);
and gate_295(n385,n139,n384);
not gate_296(n386,n385);
and gate_297(n387,n381,n386);
and gate_298(n388,n155,n270);
and gate_299(n389,pi21,n388);
and gate_300(n390,pi25,n389);
and gate_301(n391,n139,n390);
not gate_302(n392,n391);
and gate_303(n393,pi26,pi30);
and gate_304(n394,n155,n241);
and gate_305(n395,pi21,n394);
and gate_306(n396,n120,n395);
and gate_307(n397,n393,n396);
not gate_308(n398,n397);
and gate_309(n399,n392,n398);
and gate_310(n400,n387,n399);
and gate_311(n401,n107,n215);
and gate_312(n402,pi22,n350);
and gate_313(n403,n119,n402);
and gate_314(n404,n401,n403);
and gate_315(n405,n139,n404);
not gate_316(n406,n405);
and gate_317(n407,pi10,pi18);
and gate_318(n408,n111,n407);
and gate_319(n409,n352,n408);
and gate_320(n410,pi20,n409);
and gate_321(n411,pi25,n410);
and gate_322(n412,n358,n411);
not gate_323(n413,n412);
and gate_324(n414,n406,n413);
and gate_325(n415,n155,n233);
and gate_326(n416,pi21,n415);
and gate_327(n417,n120,n416);
and gate_328(n418,n393,n417);
not gate_329(n419,n418);
and gate_330(n420,n136,n318);
and gate_331(n421,n119,n420);
and gate_332(n422,n401,n421);
and gate_333(po41,n139,n422);
not gate_334(n424,po41);
and gate_335(n425,n419,n424);
and gate_336(n426,n414,n425);
and gate_337(n427,n400,n426);
and gate_338(n428,n378,n427);
and gate_339(n429,n327,n428);
not gate_340(po06,n429);
and gate_341(n431,n386,n392);
and gate_342(n432,n413,n431);
and gate_343(n433,n257,n276);
and gate_344(n434,n369,n433);
and gate_345(n435,n432,n434);
not gate_346(po07,n435);
and gate_347(n437,n247,n257);
and gate_348(n438,n230,n437);
and gate_349(n439,n269,n287);
and gate_350(n440,n323,n348);
and gate_351(n441,n439,n440);
and gate_352(n442,n438,n441);
and gate_353(n443,n398,n424);
and gate_354(n444,n387,n443);
and gate_355(n445,n356,n375);
and gate_356(n446,n414,n445);
and gate_357(n447,n444,n446);
and gate_358(n448,n442,n447);
not gate_359(po08,n448);
and gate_360(n450,n214,n340);
not gate_361(po09,n450);
and gate_362(n452,n110,n111);
and gate_363(n453,n112,n452);
and gate_364(n454,pi21,n453);
and gate_365(n455,pi22,n454);
and gate_366(n456,n119,n455);
and gate_367(n457,pi29,n456);
and gate_368(n458,pi30,n457);
not gate_369(n459,n458);
and gate_370(n460,n101,n456);
and gate_371(n461,n258,n460);
and gate_372(n462,n128,n461);
and gate_373(n463,n129,n462);
and gate_374(n464,n131,n463);
and gate_375(n465,n130,n464);
and gate_376(n466,n132,n465);
and gate_377(n467,n133,n466);
not gate_378(n468,n467);
and gate_379(n469,pi44,n467);
not gate_380(n470,n469);
and gate_381(n471,n459,n470);
and gate_382(n472,pi42,n464);
not gate_383(n473,n472);
and gate_384(n474,pi39,n462);
and gate_385(n475,n131,n474);
not gate_386(n476,n475);
and gate_387(n477,n473,n476);
and gate_388(n478,n471,n477);
and gate_389(n479,pi38,n461);
not gate_390(n480,n479);
and gate_391(n481,pi09,n456);
and gate_392(n482,n139,n481);
and gate_393(n483,n122,n482);
and gate_394(n484,n124,n483);
not gate_395(n485,n484);
and gate_396(n486,pi39,n484);
not gate_397(n487,n486);
and gate_398(n488,pi41,n462);
not gate_399(n489,n488);
and gate_400(n490,n487,n489);
and gate_401(n491,n480,n490);
and gate_402(n492,pi30,n227);
not gate_403(n493,n492);
and gate_404(n494,pi27,n218);
and gate_405(n495,n139,n494);
not gate_406(n496,n495);
and gate_407(n497,n139,n460);
not gate_408(n498,n497);
and gate_409(n499,n496,n498);
and gate_410(n500,n493,n499);
and gate_411(n501,n491,n500);
and gate_412(n502,n478,n501);
and gate_413(n503,n120,n226);
and gate_414(n504,n121,n503);
not gate_415(n505,n504);
and gate_416(n506,pi26,n252);
and gate_417(n507,pi28,n506);
and gate_418(n508,n258,n507);
not gate_419(n509,n508);
and gate_420(n510,n505,n509);
and gate_421(n511,n119,n506);
and gate_422(n512,pi29,n511);
and gate_423(n513,pi30,n512);
not gate_424(n514,n513);
and gate_425(n515,pi22,n252);
and gate_426(n516,pi29,n515);
and gate_427(n517,pi30,n516);
not gate_428(n518,n517);
and gate_429(n519,pi30,n254);
not gate_430(n520,n519);
and gate_431(n521,n518,n520);
and gate_432(n522,n514,n521);
and gate_433(n523,n510,n522);
and gate_434(n524,pi20,n135);
and gate_435(n525,n113,n524);
and gate_436(n526,pi22,n525);
and gate_437(n527,pi28,n526);
and gate_438(n528,pi29,n527);
and gate_439(n529,pi30,n528);
not gate_440(n530,n529);
and gate_441(n531,n119,n526);
and gate_442(n532,pi29,n531);
and gate_443(n533,pi30,n532);
not gate_444(n534,n533);
and gate_445(n535,n112,n135);
and gate_446(n536,pi01,n535);
and gate_447(n537,n113,n536);
and gate_448(n538,pi23,n537);
and gate_449(n539,n258,n538);
not gate_450(n540,n539);
and gate_451(n541,n534,n540);
and gate_452(n542,n530,n541);
and gate_453(po20,pi30,n295);
not gate_454(n544,po20);
and gate_455(n545,pi28,n301);
and gate_456(po21,n258,n545);
not gate_457(n547,po21);
and gate_458(n548,n544,n547);
and gate_459(n549,n306,n548);
and gate_460(n550,n542,n549);
and gate_461(n551,n523,n550);
and gate_462(n552,n502,n551);
and gate_463(n553,n113,n453);
and gate_464(n554,n119,n553);
and gate_465(n555,pi29,n554);
and gate_466(n556,pi30,n555);
not gate_467(n557,n556);
and gate_468(n558,pi20,n452);
and gate_469(n559,n113,n558);
and gate_470(n560,n119,pi29);
and gate_471(n561,n559,n560);
and gate_472(n562,pi30,n561);
not gate_473(n563,n562);
and gate_474(n564,pi28,n559);
and gate_475(n565,n258,n564);
not gate_476(n566,n565);
and gate_477(n567,n563,n566);
and gate_478(n568,pi22,n537);
and gate_479(n569,n258,n568);
not gate_480(n570,n569);
and gate_481(n571,n567,n570);
and gate_482(n572,pi28,n553);
and gate_483(n573,n258,n572);
not gate_484(n574,n573);
and gate_485(n575,n571,n574);
and gate_486(n576,n557,n575);
and gate_487(n577,n103,n290);
and gate_488(n578,pi21,n577);
and gate_489(n579,n142,n578);
and gate_490(n580,pi29,n579);
not gate_491(n581,n580);
and gate_492(n582,pi11,n350);
and gate_493(n583,n142,n582);
and gate_494(n584,pi29,n583);
not gate_495(n585,n584);
and gate_496(n586,n581,n585);
and gate_497(n587,pi25,n582);
and gate_498(n588,n560,n587);
and gate_499(n589,n121,n588);
not gate_500(n590,n589);
and gate_501(n591,pi21,n217);
and gate_502(n592,pi29,n591);
not gate_503(n593,n592);
and gate_504(n594,n121,n592);
not gate_505(n595,n594);
and gate_506(n596,n590,n595);
and gate_507(n597,n586,n596);
and gate_508(n598,n576,n597);
and gate_509(n599,pi29,n403);
and gate_510(n600,n121,n599);
not gate_511(n601,n600);
and gate_512(n602,pi25,n578);
and gate_513(n603,n560,n602);
not gate_514(n604,n603);
and gate_515(n605,n121,n603);
not gate_516(n606,n605);
and gate_517(n607,n601,n606);
and gate_518(n608,pi29,n173);
and gate_519(n609,n121,n608);
not gate_520(n610,n609);
and gate_521(n611,pi28,n136);
and gate_522(n612,pi29,n611);
not gate_523(n613,n612);
and gate_524(n614,n121,n612);
not gate_525(n615,n614);
and gate_526(n616,pi29,n421);
not gate_527(n617,n616);
and gate_528(n618,n121,n616);
not gate_529(n619,n618);
and gate_530(n620,n615,n619);
and gate_531(n621,n610,n620);
and gate_532(n622,n607,n621);
and gate_533(n623,pi21,n558);
and gate_534(n624,pi26,n623);
and gate_535(n625,pi29,n624);
not gate_536(n626,n625);
and gate_537(n627,pi30,n625);
not gate_538(n628,n627);
and gate_539(n629,pi21,n536);
and gate_540(n630,n336,n629);
and gate_541(n631,n139,n630);
not gate_542(n632,n631);
and gate_543(n633,n628,n632);
and gate_544(n634,pi24,n623);
and gate_545(n635,pi29,n634);
not gate_546(n636,n635);
and gate_547(n637,n121,n635);
not gate_548(n638,n637);
and gate_549(n639,pi22,n629);
and gate_550(n640,n119,n639);
and gate_551(n641,n139,n640);
not gate_552(n642,n641);
and gate_553(n643,n638,n642);
and gate_554(n644,n117,n623);
and gate_555(n645,pi29,n644);
not gate_556(n646,n645);
and gate_557(n647,n121,n645);
not gate_558(n648,n647);
and gate_559(n649,n121,n625);
not gate_560(n650,n649);
and gate_561(n651,n648,n650);
and gate_562(n652,n643,n651);
and gate_563(n653,n633,n652);
and gate_564(n654,n622,n653);
and gate_565(n655,n598,n654);
and gate_566(n656,n552,n655);
not gate_567(po10,n656);
and gate_568(n658,n120,n507);
and gate_569(n659,n121,n658);
not gate_570(n660,n659);
and gate_571(n661,n514,n660);
and gate_572(n662,pi28,n120);
and gate_573(n663,n302,n662);
and gate_574(n664,n121,n663);
not gate_575(n665,n664);
and gate_576(n666,n306,n665);
and gate_577(n667,n534,n666);
and gate_578(n668,n661,n667);
and gate_579(n669,pi43,n466);
and gate_580(n670,n134,n669);
not gate_581(n671,n670);
and gate_582(n672,n95,n162);
and gate_583(n673,n113,n672);
and gate_584(n674,pi27,n673);
and gate_585(n675,n120,n674);
and gate_586(n676,n121,n675);
not gate_587(n677,n676);
and gate_588(n678,n505,n677);
and gate_589(n679,n496,n678);
and gate_590(n680,n671,n679);
and gate_591(n681,n668,n680);
and gate_592(n682,n557,n574);
and gate_593(n683,n595,n682);
and gate_594(n684,n567,n683);
and gate_595(n685,pi30,n588);
not gate_596(n686,n685);
and gate_597(n687,n586,n686);
and gate_598(n688,n684,n687);
and gate_599(n689,n681,n688);
and gate_600(n690,pi30,n599);
not gate_601(n691,n690);
and gate_602(n692,pi30,n608);
not gate_603(n693,n692);
and gate_604(n694,n601,n693);
and gate_605(n695,n691,n694);
and gate_606(n696,n604,n695);
and gate_607(n697,n610,n617);
and gate_608(n698,n613,n697);
and gate_609(n699,n696,n698);
and gate_610(n700,pi21,n535);
and gate_611(n701,pi22,n700);
and gate_612(n702,n314,n701);
not gate_613(n703,n702);
and gate_614(n704,n632,n703);
and gate_615(n705,pi30,n635);
not gate_616(n706,n705);
and gate_617(n707,n642,n706);
and gate_618(n708,n336,n700);
and gate_619(n709,n258,n708);
not gate_620(n710,n709);
and gate_621(n711,n707,n710);
and gate_622(n712,n704,n711);
and gate_623(n713,n626,n646);
and gate_624(n714,n638,n713);
and gate_625(n715,n712,n714);
and gate_626(n716,n699,n715);
and gate_627(n717,n689,n716);
not gate_628(po11,n717);
and gate_629(n719,n509,n660);
and gate_630(n720,n505,n719);
and gate_631(n721,n522,n547);
and gate_632(n722,n720,n721);
and gate_633(n723,n493,n677);
and gate_634(n724,n468,n723);
and gate_635(n725,n499,n724);
and gate_636(n726,n722,n725);
and gate_637(n727,n544,n666);
and gate_638(n728,n542,n727);
and gate_639(n729,n593,n682);
and gate_640(n730,n571,n729);
and gate_641(n731,n728,n730);
and gate_642(n732,n726,n731);
and gate_643(n733,pi30,n603);
not gate_644(n734,n733);
and gate_645(n735,n590,n734);
and gate_646(n736,n686,n735);
and gate_647(n737,n606,n691);
and gate_648(n738,n694,n737);
and gate_649(n739,n736,n738);
and gate_650(n740,n235,n407);
and gate_651(n741,pi21,n740);
and gate_652(n742,pi25,n741);
and gate_653(n743,pi30,n742);
not gate_654(n744,n743);
and gate_655(n745,pi21,n251);
and gate_656(n746,n393,n745);
not gate_657(n747,n746);
and gate_658(n748,n744,n747);
and gate_659(n749,n586,n748);
and gate_660(n750,n739,n749);
and gate_661(n751,pi30,n612);
not gate_662(n752,n751);
and gate_663(n753,n615,n710);
and gate_664(n754,n752,n753);
and gate_665(n755,n697,n754);
and gate_666(n756,n636,n703);
and gate_667(n757,n713,n756);
and gate_668(n758,n755,n757);
and gate_669(n759,n750,n758);
and gate_670(n760,n732,n759);
not gate_671(po12,n760);
and gate_672(n762,pi22,n300);
and gate_673(n763,pi30,n762);
not gate_674(n764,n763);
and gate_675(n765,pi23,n300);
and gate_676(n766,pi30,n765);
not gate_677(n767,n766);
and gate_678(n768,n764,n767);
and gate_679(n769,n161,n342);
and gate_680(n770,n113,n769);
and gate_681(n771,pi22,n770);
and gate_682(n772,n192,n771);
not gate_683(n773,n772);
and gate_684(n774,n530,n773);
and gate_685(n775,pi03,n110);
and gate_686(n776,n161,n775);
and gate_687(n777,n113,n776);
and gate_688(n778,pi22,n777);
and gate_689(n779,n192,n778);
not gate_690(n780,n779);
and gate_691(n781,n774,n780);
and gate_692(n782,n768,n781);
and gate_693(n783,n139,n531);
not gate_694(n784,n783);
and gate_695(n785,n336,n525);
and gate_696(n786,n139,n785);
not gate_697(n787,n786);
and gate_698(n788,n784,n787);
and gate_699(n789,n142,n525);
and gate_700(n790,n139,n789);
not gate_701(n791,n790);
and gate_702(n792,n788,n791);
and gate_703(n793,n113,n535);
and gate_704(n794,pi23,n793);
and gate_705(n795,n139,n794);
not gate_706(n796,n795);
and gate_707(n797,n570,n796);
and gate_708(n798,n540,n797);
and gate_709(n799,n792,n798);
and gate_710(n800,n782,n799);
and gate_711(n801,n590,n632);
and gate_712(n802,n744,n801);
and gate_713(n803,pi14,n118);
and gate_714(n804,n119,n803);
and gate_715(n805,n120,n804);
and gate_716(n806,n121,n805);
not gate_717(n807,n806);
and gate_718(n808,pi13,n106);
and gate_719(n809,n118,n808);
and gate_720(n810,n357,n809);
and gate_721(n811,n120,n810);
and gate_722(n812,n121,n811);
not gate_723(n813,n812);
and gate_724(n814,n807,n813);
and gate_725(n815,n642,n814);
and gate_726(n816,n802,n815);
and gate_727(n817,n336,n559);
and gate_728(n818,n139,n817);
not gate_729(n819,n818);
and gate_730(n820,pi22,n793);
and gate_731(n821,n139,n820);
not gate_732(n822,n821);
and gate_733(n823,n819,n822);
and gate_734(n824,pi30,n592);
not gate_735(n825,n824);
and gate_736(n826,n139,n554);
not gate_737(n827,n826);
and gate_738(n828,n825,n827);
and gate_739(n829,n747,n828);
and gate_740(n830,n823,n829);
and gate_741(n831,n816,n830);
and gate_742(n832,n800,n831);
and gate_743(n833,n139,n511);
not gate_744(n834,n833);
and gate_745(n835,n660,n834);
and gate_746(n836,n113,n740);
and gate_747(n837,pi25,n836);
and gate_748(n838,n139,n837);
not gate_749(n839,n838);
and gate_750(n840,n521,n839);
and gate_751(n841,n835,n840);
and gate_752(n842,n139,n515);
not gate_753(n843,n842);
and gate_754(n844,n548,n843);
and gate_755(n845,n139,n303);
not gate_756(n846,n845);
and gate_757(n847,n139,n294);
not gate_758(n848,n847);
and gate_759(n849,n846,n848);
and gate_760(n850,n665,n849);
and gate_761(n851,n844,n850);
and gate_762(n852,n841,n851);
and gate_763(n853,n139,n220);
not gate_764(n854,n853);
and gate_765(n855,n509,n854);
and gate_766(n856,n487,n855);
and gate_767(n857,n723,n856);
and gate_768(n858,n478,n857);
and gate_769(n859,n852,n858);
and gate_770(n860,n832,n859);
not gate_771(po13,n860);
and gate_772(n862,pi40,n464);
and gate_773(n863,n132,n862);
not gate_774(n864,n863);
and gate_775(n865,n132,n475);
not gate_776(n866,n865);
and gate_777(n867,n459,n866);
and gate_778(n868,n864,n867);
and gate_779(n869,pi33,n482);
not gate_780(n870,n869);
and gate_781(n871,n677,n870);
and gate_782(n872,n490,n871);
and gate_783(n873,n868,n872);
and gate_784(n874,n493,n719);
and gate_785(n875,n521,n548);
and gate_786(n876,n874,n875);
and gate_787(n877,n873,n876);
and gate_788(n878,pi30,n616);
not gate_789(n879,n878);
and gate_790(n880,n752,n879);
and gate_791(n881,n633,n880);
and gate_792(n882,pi30,n584);
not gate_793(n883,n882);
and gate_794(n884,pi30,n580);
not gate_795(n885,n884);
and gate_796(n886,n590,n885);
and gate_797(n887,n883,n886);
and gate_798(n888,n881,n887);
and gate_799(n889,n665,n774);
and gate_800(n890,n540,n570);
and gate_801(n891,n747,n780);
and gate_802(n892,n890,n891);
and gate_803(n893,n889,n892);
and gate_804(n894,n888,n893);
and gate_805(n895,n877,n894);
not gate_806(po14,n895);
and gate_807(n897,pi05,n110);
and gate_808(n898,n95,n111);
and gate_809(n899,n897,n898);
and gate_810(n900,n112,n899);
and gate_811(n901,n113,n900);
and gate_812(n902,n314,n901);
not gate_813(n903,n902);
and gate_814(n904,n334,n903);
and gate_815(n905,n682,n904);
and gate_816(n906,pi03,n555);
and gate_817(n907,n121,n906);
not gate_818(n908,n907);
and gate_819(n909,n121,n580);
not gate_820(n910,n909);
and gate_821(n911,n121,n584);
not gate_822(n912,n911);
and gate_823(n913,n910,n912);
and gate_824(n914,n595,n913);
and gate_825(n915,n908,n914);
and gate_826(n916,n905,n915);
and gate_827(n917,pi06,n775);
and gate_828(n918,n154,n917);
and gate_829(n919,n113,n918);
and gate_830(n920,n192,n919);
not gate_831(n921,n920);
and gate_832(n922,pi06,n343);
and gate_833(n923,pi20,n922);
and gate_834(n924,n113,n923);
and gate_835(n925,n192,n924);
not gate_836(n926,n925);
and gate_837(n927,n921,n926);
and gate_838(n928,n348,n822);
and gate_839(n929,n927,n928);
and gate_840(n930,pi24,n559);
and gate_841(n931,n139,n930);
not gate_842(n932,n931);
and gate_843(n933,n567,n932);
and gate_844(n934,n929,n933);
and gate_845(n935,n916,n934);
and gate_846(n936,n590,n607);
and gate_847(n937,n199,n610);
and gate_848(n938,n172,n662);
and gate_849(n939,n121,n938);
not gate_850(n940,n939);
and gate_851(n941,n619,n940);
and gate_852(n942,n937,n941);
and gate_853(n943,n936,n942);
and gate_854(n944,n615,n632);
and gate_855(n945,n814,n944);
and gate_856(n946,n652,n945);
and gate_857(n947,n943,n946);
and gate_858(n948,n935,n947);
and gate_859(n949,pi23,n454);
and gate_860(n950,n258,n949);
and gate_861(n951,n122,n950);
and gate_862(n952,n123,n951);
and gate_863(n953,n124,n952);
not gate_864(n954,n953);
and gate_865(n955,n125,n953);
and gate_866(n956,n126,n955);
and gate_867(n957,n127,n956);
and gate_868(n958,pi37,n957);
not gate_869(n959,n958);
and gate_870(n960,pi34,n953);
not gate_871(n961,n960);
and gate_872(n962,pi35,n955);
not gate_873(n963,n962);
and gate_874(n964,n961,n963);
and gate_875(n965,n959,n964);
and gate_876(n966,pi31,n950);
not gate_877(n967,n966);
and gate_878(n968,pi32,n951);
not gate_879(n969,n968);
and gate_880(n970,n967,n969);
and gate_881(n971,n139,n949);
not gate_882(n972,n971);
and gate_883(n973,n671,n972);
and gate_884(n974,n970,n973);
and gate_885(n975,n965,n974);
and gate_886(n976,n214,n496);
and gate_887(n977,pi28,n455);
and gate_888(n978,pi30,n977);
not gate_889(n979,n978);
and gate_890(n980,n314,n494);
not gate_891(n981,n980);
and gate_892(n982,n979,n981);
and gate_893(n983,n976,n982);
and gate_894(n984,pi05,pi18);
and gate_895(n985,n161,n984);
and gate_896(n986,n113,n985);
and gate_897(n987,n118,n986);
and gate_898(n988,n560,n987);
and gate_899(n989,pi30,n988);
not gate_900(n990,n989);
and gate_901(n991,pi04,n227);
and gate_902(n992,n121,n991);
not gate_903(n993,n992);
and gate_904(n994,n505,n993);
and gate_905(n995,n990,n994);
and gate_906(n996,n493,n995);
and gate_907(n997,n983,n996);
and gate_908(n998,n975,n997);
and gate_909(n999,n514,n834);
and gate_910(n1000,n509,n999);
and gate_911(n1001,n875,n1000);
and gate_912(n1002,n306,n846);
and gate_913(n1003,n120,n527);
and gate_914(n1004,pi30,n328);
and gate_915(n1005,n1003,n1004);
not gate_916(n1006,n1005);
and gate_917(n1007,n530,n1006);
and gate_918(n1008,n1002,n1007);
and gate_919(n1009,n161,n897);
and gate_920(n1010,n113,n1009);
and gate_921(n1011,pi22,n1010);
and gate_922(n1012,n314,n1011);
not gate_923(n1013,n1012);
and gate_924(n1014,n534,n1013);
and gate_925(n1015,n890,n1014);
and gate_926(n1016,n1008,n1015);
and gate_927(n1017,n1001,n1016);
and gate_928(n1018,n998,n1017);
and gate_929(n1019,n948,n1018);
not gate_930(po15,n1019);
and gate_931(n1021,pi42,n475);
not gate_932(n1022,n1021);
and gate_933(n1023,n459,n1022);
and gate_934(n1024,n470,n1023);
and gate_935(n1025,n473,n489);
and gate_936(n1026,n866,n1025);
and gate_937(n1027,n1024,n1026);
and gate_938(n1028,n487,n498);
and gate_939(n1029,n480,n1028);
and gate_940(n1030,n214,n723);
and gate_941(n1031,n981,n1030);
and gate_942(n1032,n1029,n1031);
and gate_943(n1033,n1027,n1032);
and gate_944(n1034,n121,n221);
not gate_945(n1035,n1034);
and gate_946(n1036,n854,n1035);
and gate_947(n1037,n719,n1036);
and gate_948(n1038,n995,n1037);
and gate_949(n1039,n520,n834);
and gate_950(n1040,n839,n1039);
and gate_951(n1041,n518,n844);
and gate_952(n1042,n1040,n1041);
and gate_953(n1043,n1038,n1042);
and gate_954(n1044,n1033,n1043);
and gate_955(n1045,n590,n650);
and gate_956(n1046,n814,n1045);
and gate_957(n1047,n908,n913);
and gate_958(n1048,n1046,n1047);
and gate_959(n1049,n348,n927);
and gate_960(n1050,pi22,n559);
and gate_961(po24,n139,n1050);
not gate_962(n1052,po24);
and gate_963(n1053,n258,n930);
not gate_964(n1054,n1053);
and gate_965(n1055,n1052,n1054);
and gate_966(n1056,n904,n1055);
and gate_967(n1057,n1049,n1056);
and gate_968(n1058,n1048,n1057);
and gate_969(n1059,n780,n1013);
and gate_970(n1060,n530,n1059);
and gate_971(n1061,n787,n791);
and gate_972(n1062,n890,n1061);
and gate_973(n1063,n1060,n1062);
and gate_974(n1064,n773,n1006);
and gate_975(n1065,n764,n1064);
and gate_976(n1066,n850,n1065);
and gate_977(n1067,n1063,n1066);
and gate_978(n1068,n1058,n1067);
and gate_979(n1069,n1044,n1068);
not gate_980(po16,n1069);
and gate_981(n1071,pi36,n956);
not gate_982(n1072,n1071);
and gate_983(n1073,n959,n1072);
and gate_984(n1074,n973,n1073);
and gate_985(n1075,n134,n467);
not gate_986(n1076,n1075);
and gate_987(n1077,n979,n1076);
and gate_988(n1078,n864,n870);
and gate_989(n1079,n1077,n1078);
and gate_990(n1080,n1074,n1079);
and gate_991(n1081,n496,n981);
and gate_992(n1082,n493,n1035);
and gate_993(n1083,n1081,n1082);
and gate_994(n1084,n719,n999);
and gate_995(n1085,n520,n1084);
and gate_996(n1086,n1083,n1085);
and gate_997(n1087,n1080,n1086);
and gate_998(n1088,n768,n1002);
and gate_999(n1089,n518,n665);
and gate_1000(n1090,n548,n1089);
and gate_1001(n1091,n1088,n1090);
and gate_1002(n1092,n534,n780);
and gate_1003(n1093,n774,n1092);
and gate_1004(n1094,n787,n822);
and gate_1005(n1095,n933,n1094);
and gate_1006(n1096,n1093,n1095);
and gate_1007(n1097,n1091,n1096);
and gate_1008(n1098,n1087,n1097);
and gate_1009(n1099,pi22,n745);
and gate_1010(n1100,pi30,n1099);
not gate_1011(n1101,n1100);
and gate_1012(n1102,n883,n1101);
and gate_1013(n1103,n748,n1102);
and gate_1014(n1104,n729,n1103);
and gate_1015(n1105,pi30,n938);
not gate_1016(n1106,n1105);
and gate_1017(n1107,n885,n1106);
and gate_1018(n1108,n739,n1107);
and gate_1019(n1109,n1104,n1108);
and gate_1020(n1110,pi30,n645);
not gate_1021(n1111,n1110);
and gate_1022(n1112,n650,n1111);
and gate_1023(n1113,n648,n814);
and gate_1024(n1114,n1112,n1113);
and gate_1025(n1115,n628,n638);
and gate_1026(n1116,n707,n1115);
and gate_1027(n1117,n1114,n1116);
and gate_1028(n1118,n704,n755);
and gate_1029(n1119,n1117,n1118);
and gate_1030(n1120,n1109,n1119);
and gate_1031(n1121,n1098,n1120);
not gate_1032(po17,n1121);
and gate_1033(n1123,n964,n981);
and gate_1034(n1124,n1073,n1123);
and gate_1035(n1125,n677,n854);
and gate_1036(n1126,n496,n1125);
and gate_1037(n1127,n839,n843);
and gate_1038(n1128,n514,n1127);
and gate_1039(n1129,n1126,n1128);
and gate_1040(n1130,n1124,n1129);
and gate_1041(n1131,n306,n848);
and gate_1042(n1132,n112,n408);
and gate_1043(n1133,n113,n1132);
and gate_1044(n1134,pi25,n1133);
and gate_1045(n1135,pi30,n1134);
not gate_1046(n1136,n1135);
and gate_1047(n1137,n534,n1136);
and gate_1048(n1138,n764,n1137);
and gate_1049(n1139,n1131,n1138);
and gate_1050(n1140,n799,n1139);
and gate_1051(n1141,n1130,n1140);
and gate_1052(n1142,n566,n822);
and gate_1053(n1143,n819,n932);
and gate_1054(n1144,n563,n1143);
and gate_1055(n1145,n1142,n1144);
and gate_1056(n1146,n607,n827);
and gate_1057(n1147,n683,n1146);
and gate_1058(n1148,n1145,n1147);
and gate_1059(n1149,n632,n643);
and gate_1060(n1150,n1113,n1149);
and gate_1061(n1151,n620,n1106);
and gate_1062(n1152,n937,n1151);
and gate_1063(n1153,n1150,n1152);
and gate_1064(n1154,n1148,n1153);
and gate_1065(n1155,n1141,n1154);
not gate_1066(po18,n1155);
and gate_1067(n1157,pi33,n952);
not gate_1068(n1158,n1157);
and gate_1069(n1159,n969,n1158);
and gate_1070(n1160,n963,n1159);
and gate_1071(n1161,n671,n982);
and gate_1072(n1162,n1160,n1161);
and gate_1073(n1163,n661,n854);
and gate_1074(n1164,n679,n1163);
and gate_1075(n1165,n1162,n1164);
and gate_1076(n1166,n834,n1127);
and gate_1077(n1167,n665,n1131);
and gate_1078(n1168,n1166,n1167);
and gate_1079(n1169,n788,n1092);
and gate_1080(n1170,n767,n846);
and gate_1081(n1171,n773,n1170);
and gate_1082(n1172,n1169,n1171);
and gate_1083(n1173,n1168,n1172);
and gate_1084(n1174,n1165,n1173);
and gate_1085(n1175,n619,n944);
and gate_1086(n1176,n652,n1175);
and gate_1087(n1177,n913,n937);
and gate_1088(n1178,n607,n1177);
and gate_1089(n1179,n1176,n1178);
and gate_1090(n1180,n796,n822);
and gate_1091(n1181,n540,n1180);
and gate_1092(n1182,n567,n819);
and gate_1093(n1183,n1181,n1182);
and gate_1094(n1184,n574,n1052);
and gate_1095(n1185,n1054,n1184);
and gate_1096(n1186,n595,n827);
and gate_1097(n1187,n557,n1186);
and gate_1098(n1188,n1185,n1187);
and gate_1099(n1189,n1183,n1188);
and gate_1100(n1190,n1179,n1189);
and gate_1101(n1191,n1174,n1190);
not gate_1102(po19,n1191);
and gate_1103(n1193,n470,n864);
and gate_1104(n1194,n459,n979);
and gate_1105(n1195,n1193,n1194);
and gate_1106(n1196,n973,n1076);
and gate_1107(n1197,n1195,n1196);
and gate_1108(n1198,n970,n1158);
and gate_1109(n1199,n1073,n1198);
and gate_1110(n1200,n964,n1199);
and gate_1111(n1201,n1197,n1200);
and gate_1112(n1202,n491,n870);
and gate_1113(n1203,n477,n1202);
and gate_1114(n1204,n498,n1081);
and gate_1115(n1205,n994,n1204);
and gate_1116(n1206,n1030,n1205);
and gate_1117(n1207,n1203,n1206);
and gate_1118(n1208,n1201,n1207);
and gate_1119(n1209,n990,n1036);
and gate_1120(n1210,n1084,n1209);
and gate_1121(n1211,n102,pi18);
and gate_1122(n1212,n235,n1211);
and gate_1123(n1213,n113,n1212);
and gate_1124(n1214,pi25,n1213);
and gate_1125(n1215,n139,n1214);
not gate_1126(n1216,n1215);
and gate_1127(n1217,n839,n1216);
and gate_1128(n1218,n520,n1217);
and gate_1129(n1219,n1041,n1218);
and gate_1130(n1220,n1210,n1219);
and gate_1131(n1221,n111,n1211);
and gate_1132(n1222,n112,n1221);
and gate_1133(n1223,n113,n1222);
and gate_1134(n1224,pi25,n1223);
and gate_1135(n1225,pi30,n1224);
not gate_1136(n1226,n1225);
and gate_1137(n1227,n768,n846);
and gate_1138(n1228,n1226,n1227);
and gate_1139(n1229,n1167,n1228);
and gate_1140(n1230,n1006,n1136);
and gate_1141(n1231,n791,n1013);
and gate_1142(n1232,n1230,n1231);
and gate_1143(n1233,n1093,n1232);
and gate_1144(n1234,n1229,n1233);
and gate_1145(n1235,n1220,n1234);
and gate_1146(n1236,n1208,n1235);
and gate_1147(n1237,n154,n984);
and gate_1148(n1238,pi21,n1237);
and gate_1149(n1239,n102,n1238);
and gate_1150(n1240,pi25,n1239);
and gate_1151(n1241,n119,n1240);
and gate_1152(n1242,n139,n1241);
not gate_1153(n1243,n1242);
and gate_1154(n1244,n401,n1221);
and gate_1155(n1245,pi20,n1244);
and gate_1156(n1246,pi25,n1245);
and gate_1157(n1247,n358,n1246);
not gate_1158(n1248,n1247);
and gate_1159(n1249,n1243,n1248);
and gate_1160(n1250,n737,n1249);
and gate_1161(n1251,n736,n1250);
and gate_1162(n1252,n617,n937);
and gate_1163(n1253,n693,n940);
and gate_1164(n1254,n1106,n1253);
and gate_1165(n1255,n601,n1254);
and gate_1166(n1256,n1252,n1255);
and gate_1167(n1257,n1251,n1256);
and gate_1168(n1258,n102,n136);
and gate_1169(n1259,pi25,n1258);
and gate_1170(n1260,n119,n1259);
and gate_1171(n1261,n139,n1260);
not gate_1172(n1262,n1261);
and gate_1173(n1263,n704,n1262);
and gate_1174(n1264,n642,n1263);
and gate_1175(n1265,n754,n1264);
and gate_1176(n1266,n648,n807);
and gate_1177(n1267,n102,n110);
and gate_1178(n1268,n154,n1267);
and gate_1179(n1269,pi21,n1268);
and gate_1180(n1270,pi25,n1269);
not gate_1181(n1271,n1270);
and gate_1182(n1272,n1111,n1271);
and gate_1183(n1273,n1266,n1272);
and gate_1184(n1274,n626,n636);
and gate_1185(n1275,n1273,n1274);
and gate_1186(n1276,n1265,n1275);
and gate_1187(n1277,n1257,n1276);
and gate_1188(n1278,n827,n908);
and gate_1189(n1279,n593,n1278);
and gate_1190(n1280,n557,n904);
and gate_1191(n1281,n1279,n1280);
and gate_1192(n1282,pi21,n1212);
and gate_1193(n1283,pi25,n1282);
and gate_1194(n1284,pi30,n1283);
not gate_1195(n1285,n1284);
and gate_1196(n1286,n748,n1285);
and gate_1197(n1287,n1101,n1286);
and gate_1198(n1288,n586,n1287);
and gate_1199(n1289,n1281,n1288);
and gate_1200(n1290,n788,n928);
and gate_1201(n1291,n798,n1290);
and gate_1202(n1292,n927,n1055);
and gate_1203(n1293,n1144,n1292);
and gate_1204(n1294,n1291,n1293);
and gate_1205(n1295,n1289,n1294);
and gate_1206(n1296,n1277,n1295);
and gate_1207(n1297,n1236,n1296);
not gate_1208(po22,n1297);
and gate_1209(n1299,n650,n913);
not gate_1210(po23,n1299);
and gate_1211(n1301,n834,n854);
and gate_1212(n1302,n972,n1301);
and gate_1213(n1303,n843,n848);
and gate_1214(n1304,n1217,n1303);
and gate_1215(n1305,n1302,n1304);
and gate_1216(n1306,n113,n171);
and gate_1217(n1307,pi22,n1306);
and gate_1218(n1308,pi30,n1307);
not gate_1219(n1309,n1308);
and gate_1220(n1310,n1136,n1309);
and gate_1221(n1311,n1226,n1310);
and gate_1222(n1312,n1227,n1311);
and gate_1223(n1313,n1061,n1312);
and gate_1224(n1314,n1305,n1313);
and gate_1225(n1315,n784,n1180);
and gate_1226(n1316,n932,n1052);
not gate_1227(po43,n1316);
and gate_1228(n1318,n120,n559);
and gate_1229(n1319,n393,n1318);
not gate_1230(n1320,n1319);
and gate_1231(n1321,n819,n1320);
and gate_1232(n1322,n1316,n1321);
and gate_1233(n1323,n1315,n1322);
and gate_1234(n1324,n813,n1271);
and gate_1235(n1325,n1243,n1262);
and gate_1236(n1326,n1324,n1325);
and gate_1237(n1327,pi22,n591);
and gate_1238(n1328,pi30,n1327);
not gate_1239(n1329,n1328);
and gate_1240(n1330,n827,n1329);
and gate_1241(n1331,n1248,n1285);
and gate_1242(n1332,n1330,n1331);
and gate_1243(n1333,n1326,n1332);
and gate_1244(n1334,n1323,n1333);
and gate_1245(n1335,n1314,n1334);
not gate_1246(po25,n1335);
and gate_1247(n1337,n819,n827);
and gate_1248(n1338,n784,n854);
and gate_1249(n1339,n1337,n1338);
not gate_1250(po26,n1339);
and gate_1251(n1341,n904,n908);
and gate_1252(n1342,n1049,n1341);
and gate_1253(n1343,n990,n993);
and gate_1254(n1344,n1006,n1013);
and gate_1255(n1345,n214,n1344);
and gate_1256(n1346,n1343,n1345);
and gate_1257(n1347,n1342,n1346);
not gate_1258(po27,n1347);
and gate_1259(n1349,n1077,n1198);
and gate_1260(n1350,n954,n1349);
and gate_1261(n1351,n825,n1329);
and gate_1262(n1352,n1052,n1351);
and gate_1263(n1353,n1286,n1352);
and gate_1264(n1354,n1054,n1320);
and gate_1265(n1355,n1311,n1354);
and gate_1266(n1356,n1353,n1355);
and gate_1267(n1357,n1350,n1356);
and gate_1268(n1358,n706,n1262);
and gate_1269(n1359,n703,n1358);
and gate_1270(n1360,n628,n1272);
and gate_1271(n1361,n1359,n1360);
and gate_1272(n1362,pi08,pi16);
and gate_1273(n1363,n524,n1362);
and gate_1274(n1364,pi21,n1363);
and gate_1275(n1365,pi22,n1364);
and gate_1276(n1366,n662,n1365);
and gate_1277(n1367,n121,n1366);
not gate_1278(n1368,n1367);
and gate_1279(n1369,pi07,n108);
and gate_1280(n1370,n524,n1369);
and gate_1281(n1371,pi21,n1370);
and gate_1282(n1372,pi22,n1371);
and gate_1283(n1373,n662,n1372);
and gate_1284(n1374,n121,n1373);
not gate_1285(n1375,n1374);
and gate_1286(n1376,n1368,n1375);
and gate_1287(n1377,pi22,n1009);
and gate_1288(n1378,n358,n1377);
not gate_1289(n1379,n1378);
and gate_1290(n1380,n752,n1379);
and gate_1291(n1381,n710,n1380);
and gate_1292(n1382,n1376,n1381);
and gate_1293(n1383,n1361,n1382);
and gate_1294(n1384,n350,n1362);
and gate_1295(n1385,pi28,n1384);
not gate_1296(n1386,n1385);
and gate_1297(n1387,n350,n1369);
and gate_1298(n1388,pi28,n1387);
not gate_1299(n1389,n1388);
and gate_1300(n1390,n1386,n1389);
and gate_1301(n1391,n686,n1390);
and gate_1302(n1392,n1102,n1391);
and gate_1303(n1393,n116,n1238);
and gate_1304(n1394,n119,n1393);
and gate_1305(n1395,n139,n1394);
not gate_1306(n1396,n1395);
and gate_1307(n1397,pi05,n408);
and gate_1308(n1398,pi20,n1397);
and gate_1309(n1399,pi25,n1398);
and gate_1310(n1400,n358,n1399);
not gate_1311(n1401,n1400);
and gate_1312(n1402,n1396,n1401);
and gate_1313(n1403,n1106,n1402);
and gate_1314(n1404,n1249,n1403);
and gate_1315(n1405,n1392,n1404);
and gate_1316(n1406,n1383,n1405);
and gate_1317(n1407,n1357,n1406);
not gate_1318(po28,n1407);
and gate_1319(n1409,n317,n348);
and gate_1320(n1410,n308,n1409);
and gate_1321(n1411,n224,n263);
and gate_1322(n1412,n214,n1411);
and gate_1323(n1413,n1410,n1412);
and gate_1324(n1414,n205,n364);
and gate_1325(n1415,n340,n375);
and gate_1326(n1416,n1414,n1415);
and gate_1327(n1417,n1413,n1416);
and gate_1328(n1418,n398,n419);
and gate_1329(n1419,n189,n1418);
and gate_1330(n1420,n387,n392);
and gate_1331(n1421,n1419,n1420);
and gate_1332(n1422,n195,n424);
and gate_1333(n1423,n199,n1422);
and gate_1334(n1424,n369,n414);
and gate_1335(n1425,n1423,n1424);
and gate_1336(n1426,n1421,n1425);
and gate_1337(n1427,n1417,n1426);
not gate_1338(po29,n1427);
and gate_1339(n1429,n230,n433);
and gate_1340(n1430,n298,n323);
and gate_1341(n1431,n269,n1430);
and gate_1342(n1432,n1429,n1431);
not gate_1343(po30,n1432);
and gate_1344(n1434,n230,n248);
and gate_1345(n1435,n288,n323);
and gate_1346(n1436,n1434,n1435);
not gate_1347(po31,n1436);
and gate_1348(n1438,n104,n105);
and gate_1349(n1439,n106,n1438);
and gate_1350(n1440,n118,n1439);
and gate_1351(n1441,n357,n1440);
and gate_1352(n1442,n120,n1441);
and gate_1353(po32,n121,n1442);
not gate_1354(n1444,po32);
and gate_1355(n1445,n493,n1343);
and gate_1356(n1446,n976,n1445);
not gate_1357(po33,n1446);
and gate_1358(n1448,n470,n671);
and gate_1359(n1449,n868,n1448);
and gate_1360(n1450,n480,n485);
and gate_1361(n1451,pi31,n482);
not gate_1362(n1452,n1451);
and gate_1363(n1453,n1025,n1452);
and gate_1364(n1454,n1450,n1453);
and gate_1365(n1455,n1449,n1454);
and gate_1366(n1456,pi30,n503);
not gate_1367(n1457,n1456);
and gate_1368(n1458,n230,n1457);
and gate_1369(n1459,n870,n1458);
and gate_1370(n1460,n224,n247);
and gate_1371(n1461,n505,n1460);
and gate_1372(n1462,n1459,n1461);
and gate_1373(n1463,n240,n661);
and gate_1374(n1464,n288,n665);
and gate_1375(n1465,n1463,n1464);
and gate_1376(n1466,n1462,n1465);
and gate_1377(n1467,n1455,n1466);
and gate_1378(n1468,n195,n615);
and gate_1379(n1469,n879,n1468);
and gate_1380(n1470,n153,n1469);
and gate_1381(n1471,n691,n1253);
and gate_1382(n1472,n734,n885);
and gate_1383(n1473,n557,n1472);
and gate_1384(n1474,n1471,n1473);
and gate_1385(n1475,n1470,n1474);
and gate_1386(n1476,n120,n572);
and gate_1387(n1477,n121,n1476);
not gate_1388(n1478,n1477);
and gate_1389(n1479,n334,n1478);
and gate_1390(n1480,n563,n1479);
and gate_1391(n1481,n120,n564);
and gate_1392(n1482,n121,n1481);
not gate_1393(n1483,n1482);
and gate_1394(n1484,n348,n1483);
and gate_1395(n1485,n534,n1484);
and gate_1396(n1486,n1480,n1485);
and gate_1397(n1487,n306,n773);
and gate_1398(n1488,n121,n1003);
not gate_1399(n1489,n1488);
and gate_1400(n1490,n323,n1489);
and gate_1401(n1491,n780,n1490);
and gate_1402(n1492,n1487,n1491);
and gate_1403(n1493,n1486,n1492);
and gate_1404(n1494,n1475,n1493);
and gate_1405(n1495,n1467,n1494);
not gate_1406(po34,n1495);
and gate_1407(n1497,n972,n1022);
and gate_1408(n1498,n499,n1497);
and gate_1409(n1499,n230,n677);
and gate_1410(n1500,n1343,n1457);
and gate_1411(n1501,n1499,n1500);
and gate_1412(n1502,n1498,n1501);
and gate_1413(n1503,n248,n1036);
and gate_1414(n1504,n263,n834);
and gate_1415(n1505,n433,n839);
and gate_1416(n1506,n1504,n1505);
and gate_1417(n1507,n1503,n1506);
and gate_1418(n1508,n1502,n1507);
and gate_1419(n1509,n269,n843);
and gate_1420(n1510,n288,n1509);
and gate_1421(n1511,n773,n849);
and gate_1422(n1512,n309,n1511);
and gate_1423(n1513,n1510,n1512);
and gate_1424(n1514,n784,n796);
and gate_1425(n1515,n98,n343);
and gate_1426(n1516,pi20,n1515);
and gate_1427(n1517,n113,n1516);
and gate_1428(n1518,n192,n1517);
not gate_1429(n1519,n1518);
and gate_1430(n1520,n928,n1519);
and gate_1431(n1521,n1514,n1520);
and gate_1432(n1522,n323,n780);
and gate_1433(n1523,n530,n1522);
and gate_1434(n1524,n317,n1523);
and gate_1435(n1525,n1521,n1524);
and gate_1436(n1526,n1513,n1525);
and gate_1437(n1527,n1508,n1526);
and gate_1438(n1528,n112,n343);
and gate_1439(n1529,n113,n1528);
and gate_1440(n1530,n192,n1529);
not gate_1441(n1531,n1530);
and gate_1442(n1532,n334,n1531);
and gate_1443(n1533,n375,n1186);
and gate_1444(n1534,n1532,n1533);
and gate_1445(n1535,n98,n775);
and gate_1446(n1536,n154,n1535);
and gate_1447(n1537,n113,n1536);
and gate_1448(n1538,n192,n1537);
not gate_1449(n1539,n1538);
and gate_1450(n1540,n339,n1539);
and gate_1451(n1541,n1143,n1540);
and gate_1452(n1542,n1534,n1541);
and gate_1453(n1543,n356,n590);
and gate_1454(n1544,n413,n606);
and gate_1455(n1545,n369,n1544);
and gate_1456(n1546,n1543,n1545);
and gate_1457(n1547,n205,n363);
and gate_1458(n1548,n913,n1547);
and gate_1459(n1549,n1546,n1548);
and gate_1460(n1550,n1542,n1549);
and gate_1461(n1551,n419,n650);
and gate_1462(n1552,n189,n1551);
and gate_1463(n1553,n643,n1552);
and gate_1464(n1554,n400,n648);
and gate_1465(n1555,n1553,n1554);
and gate_1466(n1556,n406,n601);
and gate_1467(n1557,n937,n1556);
and gate_1468(n1558,n424,n619);
and gate_1469(n1559,n632,n1468);
and gate_1470(n1560,n1558,n1559);
and gate_1471(n1561,n1557,n1560);
and gate_1472(n1562,n1555,n1561);
and gate_1473(n1563,n1550,n1562);
and gate_1474(n1564,n1527,n1563);
not gate_1475(po35,n1564);
and gate_1476(n1566,n214,n1499);
and gate_1477(n1567,n1022,n1078);
and gate_1478(n1568,n1566,n1567);
and gate_1479(n1569,n263,n433);
and gate_1480(n1570,n660,n1035);
and gate_1481(n1571,n505,n1570);
and gate_1482(n1572,n1569,n1571);
and gate_1483(n1573,n1568,n1572);
and gate_1484(n1574,n298,n665);
and gate_1485(n1575,n269,n1574);
and gate_1486(n1576,n308,n1490);
and gate_1487(n1577,n1575,n1576);
and gate_1488(n1578,n339,n1483);
and gate_1489(n1579,n317,n1578);
and gate_1490(n1580,n375,n1478);
and gate_1491(n1581,n595,n912);
and gate_1492(n1582,n1580,n1581);
and gate_1493(n1583,n1579,n1582);
and gate_1494(n1584,n1577,n1583);
and gate_1495(n1585,n1573,n1584);
and gate_1496(n1586,n97,pi15);
and gate_1497(n1587,n524,n1586);
and gate_1498(n1588,pi22,n1587);
and gate_1499(n1589,n358,n1588);
not gate_1500(n1590,n1589);
and gate_1501(n1591,n620,n1590);
and gate_1502(n1592,n153,n1591);
and gate_1503(n1593,n638,n651);
and gate_1504(n1594,n106,n155);
and gate_1505(n1595,n113,n1594);
and gate_1506(n1596,n115,n1595);
and gate_1507(n1597,n118,n1596);
and gate_1508(n1598,n119,n1597);
and gate_1509(n1599,n120,n1598);
and gate_1510(n1600,n121,n1599);
not gate_1511(n1601,n1600);
and gate_1512(n1602,n120,n121);
and gate_1513(n1603,n106,n1306);
and gate_1514(n1604,n118,n1603);
and gate_1515(n1605,n119,n1604);
not gate_1516(n1606,n1605);
and gate_1517(n1607,n113,n809);
and gate_1518(n1608,n119,n1607);
not gate_1519(n1609,n1608);
and gate_1520(n1610,n1606,n1609);
not gate_1521(n1611,n1610);
and gate_1522(n1612,n1602,n1611);
not gate_1523(n1613,n1612);
and gate_1524(n1614,n1444,n1613);
and gate_1525(n1615,n1601,n1614);
and gate_1526(n1616,n1593,n1615);
and gate_1527(n1617,n1592,n1616);
and gate_1528(n1618,n735,n910);
and gate_1529(n1619,n99,n108);
and gate_1530(n1620,n350,n1619);
and gate_1531(n1621,pi28,n1620);
not gate_1532(n1622,n1621);
and gate_1533(n1623,n100,pi16);
and gate_1534(n1624,n350,n1623);
and gate_1535(n1625,pi28,n1624);
not gate_1536(n1626,n1625);
and gate_1537(n1627,n1622,n1626);
and gate_1538(n1628,n606,n1627);
and gate_1539(n1629,n1618,n1628);
and gate_1540(n1630,n601,n940);
and gate_1541(n1631,n350,n1586);
and gate_1542(n1632,n119,n1631);
and gate_1543(n1633,n139,n1632);
not gate_1544(n1634,n1633);
and gate_1545(n1635,n1630,n1634);
and gate_1546(n1636,n524,n1623);
and gate_1547(n1637,pi21,n1636);
and gate_1548(n1638,pi22,n1637);
and gate_1549(n1639,n662,n1638);
and gate_1550(n1640,n121,n1639);
not gate_1551(n1641,n1640);
and gate_1552(n1642,n524,n1619);
and gate_1553(n1643,pi21,n1642);
and gate_1554(n1644,pi22,n1643);
and gate_1555(n1645,n662,n1644);
and gate_1556(n1646,n121,n1645);
not gate_1557(n1647,n1646);
and gate_1558(n1648,n1641,n1647);
and gate_1559(n1649,n610,n1648);
and gate_1560(n1650,n1635,n1649);
and gate_1561(n1651,n1629,n1650);
and gate_1562(n1652,n1617,n1651);
and gate_1563(n1653,n1585,n1652);
not gate_1564(po36,n1653);
and gate_1565(n1655,n1196,n1198);
and gate_1566(n1656,n954,n1655);
and gate_1567(n1657,n1026,n1450);
and gate_1568(n1658,n1022,n1195);
and gate_1569(n1659,n1657,n1658);
and gate_1570(n1660,n1656,n1659);
and gate_1571(n1661,n870,n1452);
and gate_1572(n1662,n1204,n1661);
and gate_1573(n1663,n993,n1458);
and gate_1574(n1664,n1030,n1663);
and gate_1575(n1665,n1662,n1664);
and gate_1576(n1666,n224,n990);
and gate_1577(n1667,n505,n1666);
and gate_1578(n1668,n855,n1035);
and gate_1579(n1669,n1667,n1668);
and gate_1580(n1670,n248,n1504);
and gate_1581(n1671,n661,n1670);
and gate_1582(n1672,n1669,n1671);
and gate_1583(n1673,n1665,n1672);
and gate_1584(n1674,n1660,n1673);
and gate_1585(n1675,n433,n1218);
and gate_1586(n1676,n518,n547);
and gate_1587(n1677,n1510,n1676);
and gate_1588(n1678,n1675,n1677);
and gate_1589(n1679,n544,n1574);
and gate_1590(n1680,n1131,n1679);
and gate_1591(n1681,n1312,n1680);
and gate_1592(n1682,n1678,n1681);
and gate_1593(n1683,n1064,n1523);
and gate_1594(n1684,n317,n534);
and gate_1595(n1685,n1489,n1684);
and gate_1596(n1686,n1013,n1061);
and gate_1597(n1687,n1685,n1686);
and gate_1598(n1688,n1683,n1687);
and gate_1599(n1689,n1483,n1539);
and gate_1600(n1690,n1519,n1689);
and gate_1601(n1691,n1049,n1690);
and gate_1602(n1692,n1142,n1514);
and gate_1603(n1693,n890,n1692);
and gate_1604(n1694,n1691,n1693);
and gate_1605(n1695,n1688,n1694);
and gate_1606(n1696,n1682,n1695);
and gate_1607(n1697,n1674,n1696);
and gate_1608(n1698,n339,n563);
and gate_1609(n1699,n819,n1354);
and gate_1610(n1700,n1698,n1699);
and gate_1611(n1701,n932,n1184);
and gate_1612(n1702,n1479,n1531);
and gate_1613(n1703,n1701,n1702);
and gate_1614(n1704,n1700,n1703);
and gate_1615(n1705,n375,n903);
and gate_1616(n1706,n557,n1705);
and gate_1617(n1707,n828,n908);
and gate_1618(n1708,n1706,n1707);
and gate_1619(n1709,n205,n1329);
and gate_1620(n1710,n595,n1709);
and gate_1621(n1711,n1286,n1710);
and gate_1622(n1712,n1708,n1711);
and gate_1623(n1713,n1704,n1712);
and gate_1624(n1714,n363,n885);
and gate_1625(n1715,n912,n1714);
and gate_1626(n1716,n1102,n1715);
and gate_1627(n1717,n356,n686);
and gate_1628(n1718,n369,n1717);
and gate_1629(n1719,n1618,n1718);
and gate_1630(n1720,n1716,n1719);
and gate_1631(n1721,n1248,n1390);
and gate_1632(n1722,n1544,n1626);
and gate_1633(n1723,n1721,n1722);
and gate_1634(n1724,n1243,n1402);
and gate_1635(n1725,n691,n1634);
and gate_1636(n1726,n1622,n1725);
and gate_1637(n1727,n1724,n1726);
and gate_1638(n1728,n1723,n1727);
and gate_1639(n1729,n1720,n1728);
and gate_1640(n1730,n1713,n1729);
and gate_1641(n1731,n1254,n1556);
and gate_1642(n1732,n937,n1648);
and gate_1643(n1733,n1376,n1732);
and gate_1644(n1734,n1731,n1733);
and gate_1645(n1735,n710,n1468);
and gate_1646(n1736,n1263,n1735);
and gate_1647(n1737,n1380,n1590);
and gate_1648(n1738,n879,n1558);
and gate_1649(n1739,n1737,n1738);
and gate_1650(n1740,n1736,n1739);
and gate_1651(n1741,n1734,n1740);
and gate_1652(n1742,n141,n706);
and gate_1653(n1743,n642,n1742);
and gate_1654(n1744,n180,n1743);
and gate_1655(n1745,n650,n1115);
and gate_1656(n1746,n1419,n1745);
and gate_1657(n1747,n1744,n1746);
and gate_1658(n1748,n381,n646);
and gate_1659(n1749,n431,n1271);
and gate_1660(n1750,n1748,n1749);
and gate_1661(n1751,pi21,n393);
and gate_1662(n1752,n162,n1751);
not gate_1663(n1753,n1752);
and gate_1664(n1754,n807,n1753);
and gate_1665(n1755,n1615,n1754);
and gate_1666(n1756,n1750,n1755);
and gate_1667(n1757,n1747,n1756);
and gate_1668(n1758,n1741,n1757);
and gate_1669(n1759,n1730,n1758);
and gate_1670(n1760,n1697,n1759);
not gate_1671(po37,n1760);
and gate_1672(n1762,n155,n203);
not gate_1673(n1763,n1762);
and gate_1674(n1764,n113,n258);
not gate_1675(n1765,n1764);
and gate_1676(n1766,n251,n1764);
not gate_1677(n1767,n1766);
and gate_1678(n1768,n1763,n1767);
not gate_1679(n1769,n1768);
and gate_1680(n1770,n114,n116);
not gate_1681(n1771,n1770);
and gate_1682(n1772,n1769,n1771);
not gate_1683(n1773,n1772);
and gate_1684(n1774,n111,n336);
not gate_1685(n1775,n1774);
and gate_1686(n1776,pi19,pi22);
and gate_1687(n1777,pi05,n119);
not gate_1688(n1778,n1777);
and gate_1689(n1779,n1776,n1778);
not gate_1690(n1780,n1779);
and gate_1691(n1781,n1775,n1780);
not gate_1692(n1782,n1781);
and gate_1693(n1783,n110,n1782);
not gate_1694(n1784,n1783);
and gate_1695(n1785,pi19,n119);
not gate_1696(n1786,n1785);
and gate_1697(n1787,n96,n118);
and gate_1698(n1788,pi19,n1787);
not gate_1699(n1789,n1788);
and gate_1700(n1790,n143,n1789);
not gate_1701(n1791,n1790);
and gate_1702(n1792,n1786,n1791);
and gate_1703(n1793,pi18,n1792);
not gate_1704(n1794,n1793);
and gate_1705(n1795,n1784,n1794);
not gate_1706(n1796,n1795);
and gate_1707(n1797,n121,n1796);
not gate_1708(n1798,n1797);
and gate_1709(n1799,pi18,n1785);
and gate_1710(n1800,n97,n118);
and gate_1711(n1801,pi30,n1800);
and gate_1712(n1802,n1799,n1801);
not gate_1713(n1803,n1802);
and gate_1714(n1804,n1798,n1803);
not gate_1715(n1805,n1804);
and gate_1716(n1806,pi29,n1805);
not gate_1717(n1807,n1806);
and gate_1718(n1808,pi19,n209);
not gate_1719(n1809,n1808);
and gate_1720(n1810,n111,pi28);
and gate_1721(n1811,pi11,n1810);
and gate_1722(n1812,n393,n1811);
not gate_1723(n1813,n1812);
and gate_1724(n1814,n1809,n1813);
not gate_1725(n1815,n1814);
and gate_1726(n1816,pi18,n1815);
not gate_1727(n1817,n1816);
and gate_1728(n1818,n110,n1810);
and gate_1729(n1819,n1004,n1818);
not gate_1730(n1820,n1819);
and gate_1731(n1821,n1817,n1820);
not gate_1732(n1822,n1821);
and gate_1733(n1823,n120,n1822);
not gate_1734(n1824,n1823);
and gate_1735(n1825,n1807,n1824);
not gate_1736(n1826,n1825);
and gate_1737(n1827,pi20,n1826);
not gate_1738(n1828,n1827);
and gate_1739(n1829,n97,n314);
not gate_1740(n1830,n1829);
and gate_1741(n1831,n94,n192);
not gate_1742(n1832,n1831);
and gate_1743(n1833,n1830,n1832);
not gate_1744(n1834,n1833);
and gate_1745(n1835,n898,n1834);
and gate_1746(n1836,n110,n1835);
not gate_1747(n1837,n1836);
and gate_1748(n1838,n193,n315);
not gate_1749(n1839,n1838);
and gate_1750(n1840,pi26,n1839);
and gate_1751(n1841,n216,n1840);
not gate_1752(n1842,n1841);
and gate_1753(n1843,n1837,n1842);
not gate_1754(n1844,n1843);
and gate_1755(n1845,n112,n1844);
not gate_1756(n1846,n1845);
and gate_1757(n1847,n1828,n1846);
not gate_1758(n1848,n1847);
and gate_1759(n1849,n113,n1848);
not gate_1760(n1850,n1849);
and gate_1761(n1851,n119,n351);
and gate_1762(n1852,n318,n1851);
not gate_1763(n1853,n1852);
and gate_1764(n1854,n119,n1853);
not gate_1765(n1855,n1854);
and gate_1766(n1856,pi19,n1855);
not gate_1767(n1857,n1856);
and gate_1768(n1858,pi26,n154);
not gate_1769(n1859,n1858);
and gate_1770(n1860,n1857,n1859);
not gate_1771(n1861,n1860);
and gate_1772(n1862,n110,n1861);
not gate_1773(n1863,n1862);
and gate_1774(n1864,n290,n1851);
not gate_1775(n1865,n1864);
and gate_1776(n1866,n1863,n1865);
not gate_1777(n1867,n1866);
and gate_1778(n1868,n203,n1867);
not gate_1779(n1869,n1868);
and gate_1780(n1870,n1850,n1869);
and gate_1781(n1871,n1773,n1870);
not gate_1782(n1872,n1871);
and gate_1783(n1873,n92,n1872);
not gate_1784(n1874,n1873);
and gate_1785(n1875,n114,n115);
not gate_1786(n1876,n1875);
and gate_1787(n1877,n359,n1765);
not gate_1788(n1878,n1877);
and gate_1789(n1879,n1876,n1878);
and gate_1790(n1880,n535,n1879);
and gate_1791(n1881,n93,n1880);
not gate_1792(n1882,n1881);
and gate_1793(n1883,n177,n1882);
and gate_1794(n1884,n1874,n1883);
not gate_1795(po38,n1884);
and gate_1796(n1886,n509,n993);
and gate_1797(n1887,n496,n1886);
and gate_1798(n1888,n875,n1887);
and gate_1799(n1889,n540,n1344);
and gate_1800(n1890,n575,n1889);
and gate_1801(n1891,n1888,n1890);
and gate_1802(n1892,n610,n936);
and gate_1803(n1893,n914,n1892);
and gate_1804(n1894,n1176,n1893);
and gate_1805(n1895,n1891,n1894);
not gate_1806(po39,n1895);
and gate_1807(n1897,n903,n1013);
and gate_1808(n1898,n990,n1897);
and gate_1809(n1899,n908,n1379);
and gate_1810(n1900,n1402,n1899);
and gate_1811(n1901,n1898,n1900);
not gate_1812(po40,n1901);
buf gate_1813(po42,po02);
buf gate_1814(po44,po24);
endmodule
