module top(a, b, y, clk);
	input [3:0] a, b, clk;
	output wire [3:0]y;

	assign y = b;

endmodule
