// Verilog File 
module dalu (pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
pi39,pi40,pi41,pi42,pi43,pi44,pi45,pi46,pi47,pi48,
pi49,pi50,pi51,pi52,pi53,pi54,pi55,pi56,pi57,pi58,
pi59,pi60,pi61,pi62,pi63,pi64,pi65,pi66,pi67,pi68,
pi69,pi70,pi71,pi72,pi73,pi74,po00,po01,po02,po03,
po04,po05,po06,po07,po08,po09,po10,po11,po12,po13,
po14,po15);

input pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
pi39,pi40,pi41,pi42,pi43,pi44,pi45,pi46,pi47,pi48,
pi49,pi50,pi51,pi52,pi53,pi54,pi55,pi56,pi57,pi58,
pi59,pi60,pi61,pi62,pi63,pi64,pi65,pi66,pi67,pi68,
pi69,pi70,pi71,pi72,pi73,pi74;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15;

wire n91,n92,n93,n94,n95,n96,n97,n98,n99,
n100,n101,n102,n103,n104,n105,n106,n107,n108,n109,
n110,n111,n112,n113,n114,n115,n116,n117,n118,n119,
n120,n121,n122,n123,n124,n125,n126,n127,n128,n129,
n130,n131,n132,n133,n134,n135,n136,n137,n138,n139,
n140,n141,n142,n143,n144,n145,n146,n147,n148,n149,
n150,n151,n152,n153,n154,n155,n156,n157,n158,n159,
n160,n161,n162,n163,n164,n165,n166,n167,n168,n169,
n170,n171,n172,n173,n174,n175,n176,n177,n178,n179,
n180,n181,n182,n183,n184,n185,n186,n187,n188,n189,
n190,n191,n192,n193,n194,n195,n196,n197,n198,n199,
n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,
n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,
n220,n221,n222,n223,n224,n225,n226,n227,n228,n229,
n230,n231,n232,n233,n234,n235,n236,n237,n238,n239,
n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,
n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,
n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,
n270,n271,n272,n273,n274,n275,n276,n277,n278,n279,
n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,
n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,
n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,
n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,
n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,
n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,
n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,
n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,
n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,
n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,
n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,
n390,n391,n392,n393,n394,n395,n396,n397,n398,n399,
n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,
n410,n411,n412,n413,n414,n415,n416,n417,n418,n419,
n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,
n430,n431,n432,n433,n434,n435,n436,n437,n438,n439,
n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,
n450,n451,n452,n453,n454,n455,n456,n457,n458,n459,
n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,
n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,
n480,n481,n482,n483,n484,n485,n486,n487,n488,n489,
n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,
n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,
n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,
n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,
n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,
n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,
n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,
n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,
n570,n571,n572,n573,n574,n575,n576,n577,n578,n579,
n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,
n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,
n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,
n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,
n620,n621,n622,n623,n624,n625,n626,n627,n628,n629,
n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,
n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,
n650,n651,n652,n653,n654,n655,n656,n657,n658,n659,
n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,
n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,
n680,n681,n682,n683,n684,n685,n686,n687,n688,n689,
n690,n691,n692,n693,n694,n695,n696,n697,n698,n699,
n700,n701,n702,n703,n704,n705,n706,n707,n708,n709,
n710,n711,n712,n713,n714,n715,n716,n717,n718,n719,
n720,n721,n722,n723,n724,n725,n726,n727,n728,n729,
n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,
n740,n741,n742,n743,n744,n745,n746,n747,n748,n749,
n750,n751,n752,n753,n754,n755,n756,n757,n758,n759,
n760,n761,n762,n763,n764,n765,n766,n767,n768,n769,
n770,n771,n772,n773,n774,n775,n776,n777,n778,n779,
n780,n781,n782,n783,n784,n785,n786,n787,n788,n789,
n790,n791,n792,n793,n794,n795,n796,n797,n798,n799,
n800,n801,n802,n803,n804,n805,n806,n807,n808,n809,
n810,n811,n812,n813,n814,n815,n816,n817,n818,n819,
n820,n821,n822,n823,n824,n825,n826,n827,n828,n829,
n830,n831,n832,n833,n834,n835,n836,n837,n838,n839,
n840,n841,n842,n843,n844,n845,n846,n847,n848,n849,
n850,n851,n852,n853,n854,n855,n856,n857,n858,n859,
n860,n861,n862,n863,n864,n865,n866,n867,n868,n869,
n870,n871,n872,n873,n874,n875,n876,n877,n878,n879,
n880,n881,n882,n883,n884,n885,n886,n887,n888,n889,
n890,n891,n892,n893,n894,n895,n896,n897,n898,n899,
n900,n901,n902,n903,n904,n905,n906,n907,n908,n909,
n910,n911,n912,n913,n914,n915,n916,n917,n918,n919,
n920,n921,n922,n923,n924,n925,n926,n927,n928,n929,
n930,n931,n932,n933,n934,n935,n936,n937,n938,n939,
n940,n941,n942,n943,n944,n945,n946,n947,n948,n949,
n950,n951,n952,n953,n954,n955,n956,n957,n958,n959,
n960,n961,n962,n963,n964,n965,n966,n967,n968,n969,
n970,n971,n972,n973,n974,n975,n976,n977,n978,n979,
n980,n981,n982,n983,n984,n985,n986,n987,n988,n989,
n990,n991,n992,n993,n994,n995,n996,n997,n998,n999,
n1000,n1001,n1002,n1003,n1004,n1005,n1006,n1007,n1008,n1009,
n1010,n1011,n1012,n1013,n1014,n1015,n1016,n1017,n1018,n1019,
n1020,n1021,n1022,n1023,n1024,n1025,n1026,n1027,n1028,n1029,
n1030,n1031,n1032,n1033,n1034,n1035,n1036,n1037,n1038,n1039,
n1040,n1041,n1042,n1043,n1044,n1045,n1046,n1047,n1048,n1049,
n1050,n1051,n1052,n1053,n1054,n1055,n1056,n1057,n1058,n1059,
n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,n1069,
n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,n1079,
n1080,n1081,n1082,n1083,n1084,n1085,n1086,n1087,n1088,n1089,
n1090,n1091,n1092,n1093,n1094,n1095,n1096,n1097,n1098,n1099,
n1100,n1101,n1102,n1103,n1104,n1105,n1106,n1107,n1108,n1109,
n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,n1118,n1119,
n1120,n1121,n1122,n1123,n1124,n1125,n1126,n1127,n1128,n1129,
n1130,n1131,n1132,n1133,n1134,n1135,n1136,n1137,n1138,n1139,
n1140,n1141,n1142,n1143,n1144,n1145,n1146,n1147,n1148,n1149,
n1150,n1151,n1152,n1153,n1154,n1155,n1156,n1157,n1158,n1159,
n1160,n1161,n1162,n1163,n1164,n1165,n1166,n1167,n1168,n1169,
n1170,n1171,n1172,n1173,n1174,n1175,n1176,n1177,n1178,n1179,
n1180,n1181,n1182,n1183,n1184,n1185,n1186,n1187,n1188,n1189,
n1190,n1191,n1192,n1194,n1195,n1196,n1197,n1198,n1199,n1200,
n1201,n1202,n1203,n1204,n1205,n1206,n1207,n1208,n1209,n1210,
n1211,n1212,n1213,n1214,n1215,n1216,n1217,n1218,n1219,n1220,
n1221,n1222,n1223,n1224,n1225,n1226,n1227,n1228,n1229,n1230,
n1231,n1232,n1233,n1234,n1235,n1236,n1237,n1238,n1239,n1240,
n1241,n1242,n1243,n1244,n1245,n1246,n1247,n1248,n1249,n1250,
n1251,n1252,n1253,n1254,n1255,n1256,n1258,n1259,n1260,n1261,
n1262,n1263,n1264,n1265,n1266,n1267,n1268,n1269,n1270,n1271,
n1272,n1273,n1274,n1275,n1276,n1277,n1278,n1279,n1280,n1281,
n1282,n1283,n1284,n1285,n1286,n1287,n1288,n1289,n1290,n1291,
n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,n1300,n1301,
n1302,n1303,n1304,n1305,n1306,n1307,n1308,n1309,n1310,n1311,
n1312,n1313,n1314,n1315,n1316,n1317,n1318,n1319,n1320,n1321,
n1322,n1323,n1324,n1325,n1326,n1327,n1328,n1330,n1331,n1332,
n1333,n1334,n1335,n1336,n1337,n1338,n1339,n1340,n1341,n1342,
n1343,n1344,n1345,n1346,n1347,n1348,n1349,n1350,n1351,n1352,
n1353,n1354,n1355,n1356,n1357,n1358,n1359,n1360,n1361,n1362,
n1363,n1364,n1365,n1366,n1367,n1368,n1369,n1370,n1371,n1372,
n1373,n1374,n1375,n1376,n1377,n1378,n1379,n1380,n1381,n1382,
n1383,n1384,n1385,n1386,n1387,n1388,n1389,n1390,n1391,n1392,
n1393,n1394,n1395,n1396,n1397,n1398,n1399,n1400,n1401,n1402,
n1403,n1404,n1405,n1406,n1407,n1408,n1409,n1411,n1412,n1413,
n1414,n1415,n1416,n1417,n1418,n1419,n1420,n1421,n1422,n1423,
n1424,n1425,n1426,n1427,n1428,n1429,n1430,n1431,n1432,n1433,
n1434,n1435,n1436,n1437,n1438,n1439,n1440,n1441,n1442,n1443,
n1444,n1445,n1446,n1447,n1448,n1449,n1450,n1451,n1452,n1453,
n1454,n1455,n1456,n1457,n1458,n1459,n1460,n1461,n1462,n1463,
n1464,n1465,n1466,n1467,n1468,n1469,n1470,n1471,n1472,n1473,
n1474,n1475,n1476,n1477,n1478,n1479,n1480,n1481,n1482,n1483,
n1484,n1485,n1486,n1487,n1488,n1489,n1490,n1491,n1492,n1493,
n1494,n1495,n1496,n1497,n1498,n1500,n1501,n1502,n1503,n1504,
n1505,n1506,n1507,n1508,n1509,n1510,n1511,n1512,n1513,n1514,
n1515,n1516,n1517,n1518,n1519,n1520,n1521,n1522,n1523,n1524,
n1525,n1526,n1527,n1528,n1529,n1530,n1531,n1532,n1533,n1534,
n1535,n1536,n1537,n1538,n1539,n1540,n1541,n1542,n1543,n1544,
n1545,n1546,n1547,n1548,n1549,n1550,n1551,n1552,n1553,n1554,
n1555,n1556,n1557,n1558,n1559,n1560,n1561,n1562,n1563,n1564,
n1565,n1566,n1567,n1568,n1569,n1570,n1571,n1572,n1573,n1574,
n1575,n1576,n1577,n1578,n1579,n1580,n1581,n1582,n1583,n1584,
n1585,n1586,n1587,n1588,n1590,n1591,n1592,n1593,n1594,n1595,
n1596,n1597,n1598,n1599,n1600,n1601,n1602,n1603,n1604,n1605,
n1606,n1607,n1608,n1609,n1610,n1611,n1612,n1613,n1614,n1615,
n1616,n1617,n1618,n1619,n1620,n1621,n1622,n1623,n1624,n1625,
n1626,n1627,n1628,n1629,n1630,n1631,n1632,n1633,n1634,n1635,
n1636,n1637,n1638,n1639,n1640,n1641,n1642,n1643,n1644,n1645,
n1646,n1647,n1648,n1649,n1650,n1651,n1652,n1653,n1654,n1655,
n1656,n1657,n1658,n1659,n1660,n1661,n1662,n1663,n1664,n1665,
n1666,n1668,n1669,n1670,n1671,n1672,n1673,n1674,n1675,n1676,
n1677,n1678,n1679,n1680,n1681,n1682,n1683,n1684,n1685,n1686,
n1687,n1688,n1689,n1690,n1691,n1692,n1693,n1694,n1695,n1696,
n1697,n1698,n1699,n1700,n1701,n1702,n1703,n1704,n1705,n1706,
n1707,n1708,n1709,n1710,n1711,n1712,n1713,n1714,n1715,n1716,
n1717,n1718,n1719,n1720,n1721,n1722,n1723,n1724,n1725,n1726,
n1727,n1728,n1729,n1730,n1731,n1732,n1733,n1734,n1735,n1736,
n1737,n1738,n1739,n1740,n1741,n1742,n1743,n1744,n1745,n1746,
n1748,n1749,n1750,n1751,n1752,n1753,n1754,n1755,n1756,n1757,
n1758,n1759,n1760,n1761,n1762,n1763,n1764,n1765,n1766,n1767,
n1768,n1769,n1770,n1771,n1772,n1773,n1774,n1775,n1776,n1777,
n1778,n1779,n1780,n1781,n1782,n1783,n1784,n1785,n1786,n1787,
n1788,n1789,n1790,n1791,n1792,n1793,n1794,n1795,n1796,n1797,
n1798,n1799,n1800,n1801,n1802,n1803,n1804,n1805,n1806,n1807,
n1808,n1809,n1810,n1811,n1812,n1813,n1814,n1815,n1816,n1817,
n1818,n1819,n1820,n1821,n1822,n1823,n1824,n1825,n1826,n1827,
n1828,n1829,n1830,n1831,n1832,n1833,n1834,n1835,n1836,n1837,
n1838,n1840,n1841,n1842,n1843,n1844,n1845,n1846,n1847,n1848,
n1849,n1850,n1851,n1852,n1853,n1854,n1855,n1856,n1857,n1858,
n1859,n1860,n1861,n1862,n1863,n1864,n1865,n1866,n1867,n1868,
n1869,n1870,n1871,n1872,n1873,n1874,n1875,n1876,n1877,n1878,
n1879,n1880,n1881,n1882,n1883,n1884,n1885,n1886,n1887,n1888,
n1889,n1890,n1891,n1892,n1893,n1894,n1895,n1896,n1897,n1898,
n1899,n1900,n1901,n1902,n1903,n1904,n1905,n1906,n1907,n1908,
n1909,n1910,n1911,n1912,n1913,n1914,n1915,n1916,n1917,n1918,
n1920,n1921,n1922,n1923,n1924,n1925,n1926,n1927,n1928,n1929,
n1930,n1931,n1932,n1933,n1934,n1935,n1936,n1937,n1938,n1939,
n1940,n1941,n1942,n1943,n1944,n1945,n1946,n1947,n1948,n1949,
n1950,n1951,n1952,n1953,n1954,n1955,n1956,n1957,n1958,n1959,
n1960,n1961,n1962,n1963,n1964,n1965,n1966,n1967,n1968,n1969,
n1970,n1971,n1972,n1973,n1974,n1975,n1976,n1977,n1978,n1979,
n1980,n1981,n1982,n1983,n1984,n1985,n1986,n1987,n1988,n1989,
n1990,n1991,n1992,n1993,n1995,n1996,n1997,n1998,n1999,n2000,
n2001,n2002,n2003,n2004,n2005,n2006,n2007,n2008,n2009,n2010,
n2011,n2012,n2013,n2014,n2015,n2016,n2017,n2018,n2019,n2020,
n2021,n2022,n2023,n2024,n2025,n2026,n2027,n2028,n2029,n2030,
n2031,n2032,n2033,n2034,n2035,n2036,n2037,n2038,n2039,n2040,
n2041,n2042,n2043,n2044,n2045,n2046,n2047,n2048,n2049,n2050,
n2051,n2052,n2053,n2054,n2055,n2056,n2057,n2058,n2059,n2060,
n2061,n2062,n2063,n2064,n2065,n2066,n2067,n2068,n2070,n2071,
n2072,n2073,n2074,n2075,n2076,n2077,n2078,n2079,n2080,n2081,
n2082,n2083,n2084,n2085,n2086,n2087,n2088,n2089,n2090,n2091,
n2092,n2093,n2094,n2095,n2096,n2097,n2098,n2099,n2100,n2101,
n2102,n2103,n2104,n2105,n2106,n2107,n2108,n2109,n2110,n2111,
n2112,n2113,n2114,n2115,n2116,n2117,n2118,n2119,n2120,n2121,
n2122,n2123,n2124,n2125,n2126,n2127,n2128,n2129,n2130,n2131,
n2132,n2133,n2134,n2135,n2136,n2137,n2138,n2139,n2140,n2141,
n2142,n2143,n2144,n2145,n2146,n2147,n2148,n2149,n2150,n2151,
n2152,n2153,n2154,n2155,n2156,n2158,n2159,n2160,n2161,n2162,
n2163,n2164,n2165,n2166,n2167,n2168,n2169,n2170,n2171,n2172,
n2173,n2174,n2175,n2176,n2177,n2178,n2179,n2180,n2181,n2182,
n2183,n2184,n2185,n2186,n2187,n2188,n2189,n2190,n2191,n2192,
n2193,n2194,n2195,n2196,n2197,n2198,n2199,n2200,n2201,n2202,
n2203,n2204,n2205,n2206,n2207,n2208,n2209,n2210,n2211,n2212,
n2213,n2214,n2215,n2216,n2217,n2218,n2219,n2220,n2221,n2222,
n2223,n2224,n2225,n2226,n2227,n2228,n2229,n2230,n2231,n2232,
n2233,n2234,n2235,n2236,n2237,n2238,n2239,n2240,n2242,n2243,
n2244,n2245,n2246,n2247,n2248,n2249,n2250,n2251,n2252,n2253,
n2254,n2255,n2256,n2257,n2258,n2259,n2260,n2261,n2262,n2263,
n2264,n2265,n2266,n2267,n2268,n2269,n2270,n2271,n2272,n2273,
n2274,n2275,n2276,n2277,n2278,n2279,n2280,n2281,n2282,n2283,
n2284,n2285,n2286,n2287,n2288,n2289,n2290,n2291,n2292,n2293,
n2294,n2295,n2296,n2297,n2298,n2299,n2300,n2301,n2302,n2303,
n2304,n2305,n2306,n2307,n2308,n2309,n2310,n2311,n2312,n2313,
n2314,n2315,n2316,n2317,n2318,n2320,n2321,n2322,n2323,n2324,
n2325,n2326,n2327,n2328,n2329,n2330,n2331,n2332,n2333,n2334,
n2335,n2336,n2337,n2338,n2339,n2340,n2341,n2342,n2343,n2344,
n2345,n2346,n2347,n2348,n2349,n2350,n2351,n2352,n2353,n2354,
n2355,n2356,n2357,n2358,n2359,n2360,n2361,n2362,n2363,n2364,
n2365,n2366,n2367,n2368,n2369,n2370,n2371,n2372,n2373,n2374,
n2375,n2376,n2377,n2378,n2379,n2380,n2381,n2382,n2383,n2384,
n2385,n2386,n2387;
not gate_0(n91,pi64);
not gate_1(n92,pi65);
not gate_2(n93,pi66);
not gate_3(n94,pi67);
not gate_4(n95,pi68);
not gate_5(n96,pi69);
not gate_6(n97,pi70);
not gate_7(n98,pi71);
not gate_8(n99,pi72);
not gate_9(n100,pi73);
not gate_10(n101,pi74);
and gate_11(n102,n93,n94);
not gate_12(n103,n102);
and gate_13(n104,pi65,n102);
and gate_14(n105,n97,pi71);
not gate_15(n106,n105);
and gate_16(n107,pi01,n105);
not gate_17(n108,n107);
and gate_18(n109,pi33,pi70);
not gate_19(n110,n109);
and gate_20(n111,n98,n109);
not gate_21(n112,n111);
and gate_22(n113,n108,n112);
not gate_23(n114,n113);
and gate_24(n115,n96,n114);
and gate_25(n116,pi68,n115);
not gate_26(n117,n116);
and gate_27(n118,pi00,n105);
not gate_28(n119,n118);
and gate_29(n120,pi32,pi70);
not gate_30(n121,n120);
and gate_31(n122,n98,n120);
not gate_32(n123,n122);
and gate_33(n124,n119,n123);
not gate_34(n125,n124);
and gate_35(n126,n96,n125);
and gate_36(n127,pi68,n126);
not gate_37(n128,n127);
and gate_38(n129,n117,n127);
not gate_39(n130,n129);
and gate_40(n131,n116,n128);
not gate_41(n132,n131);
and gate_42(n133,n130,n132);
not gate_43(n134,n133);
and gate_44(n135,pi02,n105);
not gate_45(n136,n135);
and gate_46(n137,pi34,pi70);
not gate_47(n138,n137);
and gate_48(n139,n98,n137);
not gate_49(n140,n139);
and gate_50(n141,n136,n140);
not gate_51(n142,n141);
and gate_52(n143,n96,n142);
and gate_53(n144,pi68,n143);
not gate_54(n145,n144);
and gate_55(n146,n127,n145);
not gate_56(n147,n146);
and gate_57(n148,n128,n144);
not gate_58(n149,n148);
and gate_59(n150,n147,n149);
not gate_60(n151,n150);
and gate_61(n152,pi03,n105);
not gate_62(n153,n152);
and gate_63(n154,pi35,pi70);
not gate_64(n155,n154);
and gate_65(n156,n98,n154);
not gate_66(n157,n156);
and gate_67(n158,n153,n157);
not gate_68(n159,n158);
and gate_69(n160,n96,n159);
and gate_70(n161,pi68,n160);
not gate_71(n162,n161);
and gate_72(n163,n127,n162);
not gate_73(n164,n163);
and gate_74(n165,n128,n161);
not gate_75(n166,n165);
and gate_76(n167,n164,n166);
not gate_77(n168,n167);
and gate_78(n169,pi09,n105);
not gate_79(n170,n169);
and gate_80(n171,pi41,pi70);
not gate_81(n172,n171);
and gate_82(n173,n98,n171);
not gate_83(n174,n173);
and gate_84(n175,n170,n174);
not gate_85(n176,n175);
and gate_86(n177,n96,n176);
and gate_87(n178,pi68,n177);
not gate_88(n179,n178);
and gate_89(n180,n127,n179);
not gate_90(n181,n180);
and gate_91(n182,n128,n178);
not gate_92(n183,n182);
and gate_93(n184,n181,n183);
not gate_94(n185,n184);
and gate_95(n186,pi10,n105);
not gate_96(n187,n186);
and gate_97(n188,pi42,pi70);
not gate_98(n189,n188);
and gate_99(n190,n98,n188);
not gate_100(n191,n190);
and gate_101(n192,n187,n191);
not gate_102(n193,n192);
and gate_103(n194,n96,n193);
and gate_104(n195,pi68,n194);
not gate_105(n196,n195);
and gate_106(n197,n127,n196);
not gate_107(n198,n197);
and gate_108(n199,n128,n195);
not gate_109(n200,n199);
and gate_110(n201,n198,n200);
not gate_111(n202,n201);
and gate_112(n203,n185,n202);
and gate_113(n204,pi08,n105);
not gate_114(n205,n204);
and gate_115(n206,pi40,pi70);
not gate_116(n207,n206);
and gate_117(n208,n98,n206);
not gate_118(n209,n208);
and gate_119(n210,n205,n209);
not gate_120(n211,n210);
and gate_121(n212,n96,n211);
and gate_122(n213,pi68,n212);
not gate_123(n214,n213);
and gate_124(n215,n127,n214);
not gate_125(n216,n215);
and gate_126(n217,n128,n213);
not gate_127(n218,n217);
and gate_128(n219,n216,n218);
not gate_129(n220,n219);
and gate_130(n221,pi11,n105);
not gate_131(n222,n221);
and gate_132(n223,pi43,pi70);
not gate_133(n224,n223);
and gate_134(n225,n98,n223);
not gate_135(n226,n225);
and gate_136(n227,n222,n226);
not gate_137(n228,n227);
and gate_138(n229,n96,n228);
and gate_139(n230,pi68,n229);
not gate_140(n231,n230);
and gate_141(n232,n127,n231);
not gate_142(n233,n232);
and gate_143(n234,n128,n230);
not gate_144(n235,n234);
and gate_145(n236,n233,n235);
not gate_146(n237,n236);
and gate_147(n238,n220,n237);
and gate_148(n239,n203,n238);
and gate_149(n240,pi05,n105);
not gate_150(n241,n240);
and gate_151(n242,pi37,pi70);
not gate_152(n243,n242);
and gate_153(n244,n98,n242);
not gate_154(n245,n244);
and gate_155(n246,n241,n245);
not gate_156(n247,n246);
and gate_157(n248,n96,n247);
and gate_158(n249,pi68,n248);
not gate_159(n250,n249);
and gate_160(n251,n127,n250);
not gate_161(n252,n251);
and gate_162(n253,n128,n249);
not gate_163(n254,n253);
and gate_164(n255,n252,n254);
not gate_165(n256,n255);
and gate_166(n257,pi06,n105);
not gate_167(n258,n257);
and gate_168(n259,pi38,pi70);
not gate_169(n260,n259);
and gate_170(n261,n98,n259);
not gate_171(n262,n261);
and gate_172(n263,n258,n262);
not gate_173(n264,n263);
and gate_174(n265,n96,n264);
and gate_175(n266,pi68,n265);
not gate_176(n267,n266);
and gate_177(n268,n127,n267);
not gate_178(n269,n268);
and gate_179(n270,n128,n266);
not gate_180(n271,n270);
and gate_181(n272,n269,n271);
not gate_182(n273,n272);
and gate_183(n274,n256,n273);
and gate_184(n275,pi04,n105);
not gate_185(n276,n275);
and gate_186(n277,pi36,pi70);
not gate_187(n278,n277);
and gate_188(n279,n98,n277);
not gate_189(n280,n279);
and gate_190(n281,n276,n280);
not gate_191(n282,n281);
and gate_192(n283,n96,n282);
and gate_193(n284,pi68,n283);
not gate_194(n285,n284);
and gate_195(n286,n127,n285);
not gate_196(n287,n286);
and gate_197(n288,n128,n284);
not gate_198(n289,n288);
and gate_199(n290,n287,n289);
not gate_200(n291,n290);
and gate_201(n292,pi07,n105);
not gate_202(n293,n292);
and gate_203(n294,pi39,pi70);
not gate_204(n295,n294);
and gate_205(n296,n98,n294);
not gate_206(n297,n296);
and gate_207(n298,n293,n297);
not gate_208(n299,n298);
and gate_209(n300,n96,n299);
and gate_210(n301,pi68,n300);
not gate_211(n302,n301);
and gate_212(n303,n127,n302);
not gate_213(n304,n303);
and gate_214(n305,n128,n301);
not gate_215(n306,n305);
and gate_216(n307,n304,n306);
not gate_217(n308,n307);
and gate_218(n309,n291,n308);
and gate_219(n310,n274,n309);
and gate_220(n311,pi12,n105);
not gate_221(n312,n311);
and gate_222(n313,pi44,pi70);
not gate_223(n314,n313);
and gate_224(n315,n98,n313);
not gate_225(n316,n315);
and gate_226(n317,n312,n316);
not gate_227(n318,n317);
and gate_228(n319,n96,n318);
and gate_229(n320,pi68,n319);
not gate_230(n321,n320);
and gate_231(n322,n127,n321);
not gate_232(n323,n322);
and gate_233(n324,n128,n320);
not gate_234(n325,n324);
and gate_235(n326,n323,n325);
not gate_236(n327,n326);
and gate_237(n328,pi15,n105);
not gate_238(n329,n328);
and gate_239(n330,pi47,pi70);
not gate_240(n331,n330);
and gate_241(n332,n98,n330);
not gate_242(n333,n332);
and gate_243(n334,n329,n333);
not gate_244(n335,n334);
and gate_245(n336,n96,n335);
and gate_246(n337,pi68,n336);
not gate_247(n338,n337);
and gate_248(n339,n127,n338);
not gate_249(n340,n339);
and gate_250(n341,pi13,n105);
not gate_251(n342,n341);
and gate_252(n343,pi45,pi70);
not gate_253(n344,n343);
and gate_254(n345,n98,n343);
not gate_255(n346,n345);
and gate_256(n347,n342,n346);
not gate_257(n348,n347);
and gate_258(n349,n96,n348);
and gate_259(n350,pi68,n349);
not gate_260(n351,n350);
and gate_261(n352,n127,n351);
not gate_262(n353,n352);
and gate_263(n354,n128,n350);
not gate_264(n355,n354);
and gate_265(n356,n353,n355);
not gate_266(n357,n356);
and gate_267(n358,pi14,n105);
not gate_268(n359,n358);
and gate_269(n360,pi46,pi70);
not gate_270(n361,n360);
and gate_271(n362,n98,n360);
not gate_272(n363,n362);
and gate_273(n364,n359,n363);
not gate_274(n365,n364);
and gate_275(n366,n96,n365);
and gate_276(n367,pi68,n366);
not gate_277(n368,n367);
and gate_278(n369,n127,n368);
not gate_279(n370,n369);
and gate_280(n371,n128,n367);
not gate_281(n372,n371);
and gate_282(n373,n370,n372);
not gate_283(n374,n373);
and gate_284(n375,n357,n374);
and gate_285(n376,n339,n375);
not gate_286(n377,n376);
and gate_287(n378,n327,n376);
not gate_288(n379,n378);
and gate_289(n380,n310,n378);
not gate_290(n381,n380);
and gate_291(n382,n239,n380);
not gate_292(n383,n382);
and gate_293(n384,n168,n382);
not gate_294(n385,n384);
and gate_295(n386,n151,n384);
not gate_296(n387,n386);
and gate_297(n388,n134,n386);
not gate_298(n389,n388);
and gate_299(n390,n104,n388);
not gate_300(n391,n390);
and gate_301(n392,n97,n98);
and gate_302(n393,n96,n392);
and gate_303(n394,pi48,pi68);
and gate_304(n395,n393,n394);
not gate_305(n396,n395);
and gate_306(n397,pi48,pi70);
and gate_307(n398,pi71,n397);
not gate_308(n399,n398);
and gate_309(n400,pi70,n98);
not gate_310(n401,n400);
and gate_311(n402,n106,n401);
not gate_312(n403,n402);
and gate_313(n404,pi16,n403);
not gate_314(n405,n404);
and gate_315(n406,n399,n405);
not gate_316(n407,n406);
and gate_317(n408,n95,pi69);
and gate_318(n409,n407,n408);
not gate_319(n410,n409);
and gate_320(n411,n396,n410);
not gate_321(n412,n411);
and gate_322(n413,pi65,n412);
not gate_323(n414,n413);
and gate_324(n415,n92,n388);
not gate_325(n416,n415);
and gate_326(n417,n414,n416);
not gate_327(n418,n417);
and gate_328(n419,n103,n418);
not gate_329(n420,n419);
and gate_330(n421,n391,n420);
not gate_331(n422,n421);
and gate_332(n423,n91,n422);
not gate_333(n424,n423);
and gate_334(n425,pi64,n92);
not gate_335(n426,n425);
and gate_336(n427,n102,n412);
not gate_337(n428,n427);
and gate_338(n429,pi00,n97);
not gate_339(n430,n429);
and gate_340(n431,n121,n430);
not gate_341(n432,n431);
and gate_342(n433,n96,n432);
and gate_343(n434,pi71,n433);
not gate_344(n435,n434);
and gate_345(n436,pi69,n97);
and gate_346(n437,pi48,n436);
not gate_347(n438,n437);
and gate_348(n439,n96,pi70);
and gate_349(n440,pi16,n439);
not gate_350(n441,n440);
and gate_351(n442,n438,n441);
not gate_352(n443,n442);
and gate_353(n444,n98,n443);
not gate_354(n445,n444);
and gate_355(n446,n435,n445);
not gate_356(n447,n446);
and gate_357(n448,n95,n447);
not gate_358(n449,n448);
and gate_359(n450,pi32,pi68);
and gate_360(n451,n393,n450);
not gate_361(n452,n451);
and gate_362(n453,pi71,n120);
not gate_363(n454,n453);
and gate_364(n455,pi00,n403);
not gate_365(n456,n455);
and gate_366(n457,n454,n456);
not gate_367(n458,n457);
and gate_368(n459,n408,n458);
not gate_369(n460,n459);
and gate_370(n461,n452,n460);
not gate_371(n462,n461);
and gate_372(n463,n91,pi66);
not gate_373(n464,n463);
and gate_374(n465,n464,n426);
not gate_375(n466,n465);
and gate_376(n467,n92,pi66);
not gate_377(n468,n467);
and gate_378(n469,n94,n468);
and gate_379(n470,n466,n469);
not gate_380(n471,n470);
and gate_381(n472,n461,n470);
not gate_382(n473,n472);
and gate_383(n474,n462,n471);
not gate_384(n475,n474);
and gate_385(n476,n473,n475);
not gate_386(n477,n476);
and gate_387(n478,n449,n477);
not gate_388(n479,n478);
and gate_389(n480,n448,n476);
not gate_390(n481,n480);
and gate_391(n482,n479,n481);
not gate_392(n483,n482);
and gate_393(n484,pi33,pi68);
and gate_394(n485,n393,n484);
not gate_395(n486,n485);
and gate_396(n487,pi71,n109);
not gate_397(n488,n487);
and gate_398(n489,pi01,n403);
not gate_399(n490,n489);
and gate_400(n491,n488,n490);
not gate_401(n492,n491);
and gate_402(n493,n408,n492);
not gate_403(n494,n493);
and gate_404(n495,n486,n494);
not gate_405(n496,n495);
and gate_406(n497,n470,n495);
not gate_407(n498,n497);
and gate_408(n499,n471,n496);
not gate_409(n500,n499);
and gate_410(n501,n498,n500);
not gate_411(n502,n501);
and gate_412(n503,pi01,n97);
not gate_413(n504,n503);
and gate_414(n505,n110,n504);
not gate_415(n506,n505);
and gate_416(n507,n96,n506);
and gate_417(n508,pi71,n507);
not gate_418(n509,n508);
and gate_419(n510,pi49,n436);
not gate_420(n511,n510);
and gate_421(n512,pi17,n439);
not gate_422(n513,n512);
and gate_423(n514,n511,n513);
not gate_424(n515,n514);
and gate_425(n516,n98,n515);
not gate_426(n517,n516);
and gate_427(n518,n509,n517);
not gate_428(n519,n518);
and gate_429(n520,n95,n519);
not gate_430(n521,n520);
and gate_431(n522,n502,n520);
not gate_432(n523,n522);
and gate_433(n524,n501,n521);
not gate_434(n525,n524);
and gate_435(n526,pi34,pi68);
and gate_436(n527,n393,n526);
not gate_437(n528,n527);
and gate_438(n529,pi71,n137);
not gate_439(n530,n529);
and gate_440(n531,pi02,n403);
not gate_441(n532,n531);
and gate_442(n533,n530,n532);
not gate_443(n534,n533);
and gate_444(n535,n408,n534);
not gate_445(n536,n535);
and gate_446(n537,n528,n536);
not gate_447(n538,n537);
and gate_448(n539,n470,n537);
not gate_449(n540,n539);
and gate_450(n541,n471,n538);
not gate_451(n542,n541);
and gate_452(n543,n540,n542);
not gate_453(n544,n543);
and gate_454(n545,pi02,n97);
not gate_455(n546,n545);
and gate_456(n547,n138,n546);
not gate_457(n548,n547);
and gate_458(n549,n96,n548);
and gate_459(n550,pi71,n549);
not gate_460(n551,n550);
and gate_461(n552,pi50,n436);
not gate_462(n553,n552);
and gate_463(n554,pi18,n439);
not gate_464(n555,n554);
and gate_465(n556,n553,n555);
not gate_466(n557,n556);
and gate_467(n558,n98,n557);
not gate_468(n559,n558);
and gate_469(n560,n551,n559);
not gate_470(n561,n560);
and gate_471(n562,n95,n561);
not gate_472(n563,n562);
and gate_473(n564,n544,n562);
not gate_474(n565,n564);
and gate_475(n566,n543,n563);
not gate_476(n567,n566);
and gate_477(n568,pi35,pi68);
and gate_478(n569,n393,n568);
not gate_479(n570,n569);
and gate_480(n571,pi71,n154);
not gate_481(n572,n571);
and gate_482(n573,pi03,n403);
not gate_483(n574,n573);
and gate_484(n575,n572,n574);
not gate_485(n576,n575);
and gate_486(n577,n408,n576);
not gate_487(n578,n577);
and gate_488(n579,n570,n578);
not gate_489(n580,n579);
and gate_490(n581,n470,n579);
not gate_491(n582,n581);
and gate_492(n583,n471,n580);
not gate_493(n584,n583);
and gate_494(n585,n582,n584);
not gate_495(n586,n585);
and gate_496(n587,pi03,n97);
not gate_497(n588,n587);
and gate_498(n589,n155,n588);
not gate_499(n590,n589);
and gate_500(n591,n96,n590);
and gate_501(n592,pi71,n591);
not gate_502(n593,n592);
and gate_503(n594,pi51,n436);
not gate_504(n595,n594);
and gate_505(n596,pi19,n439);
not gate_506(n597,n596);
and gate_507(n598,n595,n597);
not gate_508(n599,n598);
and gate_509(n600,n98,n599);
not gate_510(n601,n600);
and gate_511(n602,n593,n601);
not gate_512(n603,n602);
and gate_513(n604,n95,n603);
not gate_514(n605,n604);
and gate_515(n606,n586,n604);
not gate_516(n607,n606);
and gate_517(n608,pi04,n97);
not gate_518(n609,n608);
and gate_519(n610,n278,n609);
not gate_520(n611,n610);
and gate_521(n612,n96,n611);
and gate_522(n613,pi71,n612);
not gate_523(n614,n613);
and gate_524(n615,pi52,n436);
not gate_525(n616,n615);
and gate_526(n617,pi20,n439);
not gate_527(n618,n617);
and gate_528(n619,n616,n618);
not gate_529(n620,n619);
and gate_530(n621,n98,n620);
not gate_531(n622,n621);
and gate_532(n623,n614,n622);
not gate_533(n624,n623);
and gate_534(n625,n95,n624);
not gate_535(n626,n625);
and gate_536(n627,pi36,pi68);
and gate_537(n628,n393,n627);
not gate_538(n629,n628);
and gate_539(n630,pi71,n277);
not gate_540(n631,n630);
and gate_541(n632,pi04,n403);
not gate_542(n633,n632);
and gate_543(n634,n631,n633);
not gate_544(n635,n634);
and gate_545(n636,n408,n635);
not gate_546(n637,n636);
and gate_547(n638,n629,n637);
not gate_548(n639,n638);
and gate_549(n640,n470,n638);
not gate_550(n641,n640);
and gate_551(n642,n471,n639);
not gate_552(n643,n642);
and gate_553(n644,n641,n643);
not gate_554(n645,n644);
and gate_555(n646,n625,n645);
not gate_556(n647,n646);
and gate_557(n648,n626,n644);
not gate_558(n649,n648);
and gate_559(n650,pi05,n97);
not gate_560(n651,n650);
and gate_561(n652,n243,n651);
not gate_562(n653,n652);
and gate_563(n654,n96,n653);
and gate_564(n655,pi71,n654);
not gate_565(n656,n655);
and gate_566(n657,pi53,n436);
not gate_567(n658,n657);
and gate_568(n659,pi21,n439);
not gate_569(n660,n659);
and gate_570(n661,n658,n660);
not gate_571(n662,n661);
and gate_572(n663,n98,n662);
not gate_573(n664,n663);
and gate_574(n665,n656,n664);
not gate_575(n666,n665);
and gate_576(n667,n95,n666);
not gate_577(n668,n667);
and gate_578(n669,pi37,pi68);
and gate_579(n670,n393,n669);
not gate_580(n671,n670);
and gate_581(n672,pi71,n242);
not gate_582(n673,n672);
and gate_583(n674,pi05,n403);
not gate_584(n675,n674);
and gate_585(n676,n673,n675);
not gate_586(n677,n676);
and gate_587(n678,n408,n677);
not gate_588(n679,n678);
and gate_589(n680,n671,n679);
not gate_590(n681,n680);
and gate_591(n682,n470,n680);
not gate_592(n683,n682);
and gate_593(n684,n471,n681);
not gate_594(n685,n684);
and gate_595(n686,n683,n685);
not gate_596(n687,n686);
and gate_597(n688,n668,n686);
not gate_598(n689,n688);
and gate_599(n690,n649,n689);
and gate_600(n691,pi06,n97);
not gate_601(n692,n691);
and gate_602(n693,n260,n692);
not gate_603(n694,n693);
and gate_604(n695,n96,n694);
and gate_605(n696,pi71,n695);
not gate_606(n697,n696);
and gate_607(n698,pi54,n436);
not gate_608(n699,n698);
and gate_609(n700,pi22,n439);
not gate_610(n701,n700);
and gate_611(n702,n699,n701);
not gate_612(n703,n702);
and gate_613(n704,n98,n703);
not gate_614(n705,n704);
and gate_615(n706,n697,n705);
not gate_616(n707,n706);
and gate_617(n708,n95,n707);
not gate_618(n709,n708);
and gate_619(n710,pi38,pi68);
and gate_620(n711,n393,n710);
not gate_621(n712,n711);
and gate_622(n713,pi71,n259);
not gate_623(n714,n713);
and gate_624(n715,pi06,n403);
not gate_625(n716,n715);
and gate_626(n717,n714,n716);
not gate_627(n718,n717);
and gate_628(n719,n408,n718);
not gate_629(n720,n719);
and gate_630(n721,n712,n720);
not gate_631(n722,n721);
and gate_632(n723,n470,n721);
not gate_633(n724,n723);
and gate_634(n725,n471,n722);
not gate_635(n726,n725);
and gate_636(n727,n724,n726);
not gate_637(n728,n727);
and gate_638(n729,n709,n727);
not gate_639(n730,n729);
and gate_640(n731,pi07,n97);
not gate_641(n732,n731);
and gate_642(n733,n295,n732);
not gate_643(n734,n733);
and gate_644(n735,n96,n734);
and gate_645(n736,pi71,n735);
not gate_646(n737,n736);
and gate_647(n738,pi55,n436);
not gate_648(n739,n738);
and gate_649(n740,pi23,n439);
not gate_650(n741,n740);
and gate_651(n742,n739,n741);
not gate_652(n743,n742);
and gate_653(n744,n98,n743);
not gate_654(n745,n744);
and gate_655(n746,n737,n745);
not gate_656(n747,n746);
and gate_657(n748,n95,n747);
not gate_658(n749,n748);
and gate_659(n750,pi39,pi68);
and gate_660(n751,n393,n750);
not gate_661(n752,n751);
and gate_662(n753,pi71,n294);
not gate_663(n754,n753);
and gate_664(n755,pi07,n403);
not gate_665(n756,n755);
and gate_666(n757,n754,n756);
not gate_667(n758,n757);
and gate_668(n759,n408,n758);
not gate_669(n760,n759);
and gate_670(n761,n752,n760);
not gate_671(n762,n761);
and gate_672(n763,n470,n761);
not gate_673(n764,n763);
and gate_674(n765,n471,n762);
not gate_675(n766,n765);
and gate_676(n767,n764,n766);
not gate_677(n768,n767);
and gate_678(n769,n748,n768);
not gate_679(n770,n769);
and gate_680(n771,n730,n769);
not gate_681(n772,n771);
and gate_682(n773,n708,n728);
not gate_683(n774,n773);
and gate_684(n775,n772,n774);
and gate_685(n776,n667,n687);
not gate_686(n777,n776);
and gate_687(n778,n775,n777);
not gate_688(n779,n778);
and gate_689(n780,n690,n779);
not gate_690(n781,n780);
and gate_691(n782,n647,n781);
and gate_692(n783,pi08,n97);
not gate_693(n784,n783);
and gate_694(n785,n207,n784);
not gate_695(n786,n785);
and gate_696(n787,n96,n786);
and gate_697(n788,pi71,n787);
not gate_698(n789,n788);
and gate_699(n790,pi56,n436);
not gate_700(n791,n790);
and gate_701(n792,pi24,n439);
not gate_702(n793,n792);
and gate_703(n794,n791,n793);
not gate_704(n795,n794);
and gate_705(n796,n98,n795);
not gate_706(n797,n796);
and gate_707(n798,n789,n797);
not gate_708(n799,n798);
and gate_709(n800,n95,n799);
not gate_710(n801,n800);
and gate_711(n802,pi40,pi68);
and gate_712(n803,n393,n802);
not gate_713(n804,n803);
and gate_714(n805,pi71,n206);
not gate_715(n806,n805);
and gate_716(n807,pi08,n403);
not gate_717(n808,n807);
and gate_718(n809,n806,n808);
not gate_719(n810,n809);
and gate_720(n811,n408,n810);
not gate_721(n812,n811);
and gate_722(n813,n804,n812);
not gate_723(n814,n813);
and gate_724(n815,n470,n813);
not gate_725(n816,n815);
and gate_726(n817,n471,n814);
not gate_727(n818,n817);
and gate_728(n819,n816,n818);
not gate_729(n820,n819);
and gate_730(n821,n800,n820);
not gate_731(n822,n821);
and gate_732(n823,n801,n819);
not gate_733(n824,n823);
and gate_734(n825,pi09,n97);
not gate_735(n826,n825);
and gate_736(n827,n172,n826);
not gate_737(n828,n827);
and gate_738(n829,n96,n828);
and gate_739(n830,pi71,n829);
not gate_740(n831,n830);
and gate_741(n832,pi57,n436);
not gate_742(n833,n832);
and gate_743(n834,pi25,n439);
not gate_744(n835,n834);
and gate_745(n836,n833,n835);
not gate_746(n837,n836);
and gate_747(n838,n98,n837);
not gate_748(n839,n838);
and gate_749(n840,n831,n839);
not gate_750(n841,n840);
and gate_751(n842,n95,n841);
not gate_752(n843,n842);
and gate_753(n844,pi41,pi68);
and gate_754(n845,n393,n844);
not gate_755(n846,n845);
and gate_756(n847,pi71,n171);
not gate_757(n848,n847);
and gate_758(n849,pi09,n403);
not gate_759(n850,n849);
and gate_760(n851,n848,n850);
not gate_761(n852,n851);
and gate_762(n853,n408,n852);
not gate_763(n854,n853);
and gate_764(n855,n846,n854);
not gate_765(n856,n855);
and gate_766(n857,n470,n855);
not gate_767(n858,n857);
and gate_768(n859,n471,n856);
not gate_769(n860,n859);
and gate_770(n861,n858,n860);
not gate_771(n862,n861);
and gate_772(n863,n843,n861);
not gate_773(n864,n863);
and gate_774(n865,n824,n864);
and gate_775(n866,pi10,n97);
not gate_776(n867,n866);
and gate_777(n868,n189,n867);
not gate_778(n869,n868);
and gate_779(n870,n96,n869);
and gate_780(n871,pi71,n870);
not gate_781(n872,n871);
and gate_782(n873,pi58,n436);
not gate_783(n874,n873);
and gate_784(n875,pi26,n439);
not gate_785(n876,n875);
and gate_786(n877,n874,n876);
not gate_787(n878,n877);
and gate_788(n879,n98,n878);
not gate_789(n880,n879);
and gate_790(n881,n872,n880);
not gate_791(n882,n881);
and gate_792(n883,n95,n882);
not gate_793(n884,n883);
and gate_794(n885,pi42,pi68);
and gate_795(n886,n393,n885);
not gate_796(n887,n886);
and gate_797(n888,pi71,n188);
not gate_798(n889,n888);
and gate_799(n890,pi10,n403);
not gate_800(n891,n890);
and gate_801(n892,n889,n891);
not gate_802(n893,n892);
and gate_803(n894,n408,n893);
not gate_804(n895,n894);
and gate_805(n896,n887,n895);
not gate_806(n897,n896);
and gate_807(n898,n470,n896);
not gate_808(n899,n898);
and gate_809(n900,n471,n897);
not gate_810(n901,n900);
and gate_811(n902,n899,n901);
not gate_812(n903,n902);
and gate_813(n904,n883,n903);
not gate_814(n905,n904);
and gate_815(n906,n884,n902);
not gate_816(n907,n906);
and gate_817(n908,pi11,n97);
not gate_818(n909,n908);
and gate_819(n910,n224,n909);
not gate_820(n911,n910);
and gate_821(n912,n96,n911);
and gate_822(n913,pi71,n912);
not gate_823(n914,n913);
and gate_824(n915,pi59,n436);
not gate_825(n916,n915);
and gate_826(n917,pi27,n439);
not gate_827(n918,n917);
and gate_828(n919,n916,n918);
not gate_829(n920,n919);
and gate_830(n921,n98,n920);
not gate_831(n922,n921);
and gate_832(n923,n914,n922);
not gate_833(n924,n923);
and gate_834(n925,n95,n924);
not gate_835(n926,n925);
and gate_836(n927,pi43,pi68);
and gate_837(n928,n393,n927);
not gate_838(n929,n928);
and gate_839(n930,pi71,n223);
not gate_840(n931,n930);
and gate_841(n932,pi11,n403);
not gate_842(n933,n932);
and gate_843(n934,n931,n933);
not gate_844(n935,n934);
and gate_845(n936,n408,n935);
not gate_846(n937,n936);
and gate_847(n938,n929,n937);
not gate_848(n939,n938);
and gate_849(n940,n470,n938);
not gate_850(n941,n940);
and gate_851(n942,n471,n939);
not gate_852(n943,n942);
and gate_853(n944,n941,n943);
not gate_854(n945,n944);
and gate_855(n946,n925,n945);
not gate_856(n947,n946);
and gate_857(n948,n907,n946);
not gate_858(n949,n948);
and gate_859(n950,n905,n949);
and gate_860(n951,n842,n862);
not gate_861(n952,n951);
and gate_862(n953,n950,n952);
not gate_863(n954,n953);
and gate_864(n955,n865,n954);
not gate_865(n956,n955);
and gate_866(n957,n822,n956);
and gate_867(n958,pi12,n97);
not gate_868(n959,n958);
and gate_869(n960,n314,n959);
not gate_870(n961,n960);
and gate_871(n962,n96,n961);
and gate_872(n963,pi71,n962);
not gate_873(n964,n963);
and gate_874(n965,pi60,n436);
not gate_875(n966,n965);
and gate_876(n967,pi28,n439);
not gate_877(n968,n967);
and gate_878(n969,n966,n968);
not gate_879(n970,n969);
and gate_880(n971,n98,n970);
not gate_881(n972,n971);
and gate_882(n973,n964,n972);
not gate_883(n974,n973);
and gate_884(n975,n95,n974);
not gate_885(n976,n975);
and gate_886(n977,pi44,pi68);
and gate_887(n978,n393,n977);
not gate_888(n979,n978);
and gate_889(n980,pi71,n313);
not gate_890(n981,n980);
and gate_891(n982,pi12,n403);
not gate_892(n983,n982);
and gate_893(n984,n981,n983);
not gate_894(n985,n984);
and gate_895(n986,n408,n985);
not gate_896(n987,n986);
and gate_897(n988,n979,n987);
not gate_898(n989,n988);
and gate_899(n990,n470,n988);
not gate_900(n991,n990);
and gate_901(n992,n471,n989);
not gate_902(n993,n992);
and gate_903(n994,n991,n993);
not gate_904(n995,n994);
and gate_905(n996,n975,n995);
not gate_906(n997,n996);
and gate_907(n998,n976,n994);
not gate_908(n999,n998);
and gate_909(n1000,pi13,n97);
not gate_910(n1001,n1000);
and gate_911(n1002,n344,n1001);
not gate_912(n1003,n1002);
and gate_913(n1004,n96,n1003);
and gate_914(n1005,pi71,n1004);
not gate_915(n1006,n1005);
and gate_916(n1007,pi61,n436);
not gate_917(n1008,n1007);
and gate_918(n1009,pi29,n439);
not gate_919(n1010,n1009);
and gate_920(n1011,n1008,n1010);
not gate_921(n1012,n1011);
and gate_922(n1013,n98,n1012);
not gate_923(n1014,n1013);
and gate_924(n1015,n1006,n1014);
not gate_925(n1016,n1015);
and gate_926(n1017,n95,n1016);
not gate_927(n1018,n1017);
and gate_928(n1019,pi45,pi68);
and gate_929(n1020,n393,n1019);
not gate_930(n1021,n1020);
and gate_931(n1022,pi71,n343);
not gate_932(n1023,n1022);
and gate_933(n1024,pi13,n403);
not gate_934(n1025,n1024);
and gate_935(n1026,n1023,n1025);
not gate_936(n1027,n1026);
and gate_937(n1028,n408,n1027);
not gate_938(n1029,n1028);
and gate_939(n1030,n1021,n1029);
not gate_940(n1031,n1030);
and gate_941(n1032,n470,n1030);
not gate_942(n1033,n1032);
and gate_943(n1034,n471,n1031);
not gate_944(n1035,n1034);
and gate_945(n1036,n1033,n1035);
not gate_946(n1037,n1036);
and gate_947(n1038,n1018,n1036);
not gate_948(n1039,n1038);
and gate_949(n1040,n999,n1039);
and gate_950(n1041,pi14,n97);
not gate_951(n1042,n1041);
and gate_952(n1043,n361,n1042);
not gate_953(n1044,n1043);
and gate_954(n1045,n96,n1044);
and gate_955(n1046,pi71,n1045);
not gate_956(n1047,n1046);
and gate_957(n1048,pi62,n436);
not gate_958(n1049,n1048);
and gate_959(n1050,pi30,n439);
not gate_960(n1051,n1050);
and gate_961(n1052,n1049,n1051);
not gate_962(n1053,n1052);
and gate_963(n1054,n98,n1053);
not gate_964(n1055,n1054);
and gate_965(n1056,n1047,n1055);
not gate_966(n1057,n1056);
and gate_967(n1058,n95,n1057);
not gate_968(n1059,n1058);
and gate_969(n1060,pi46,pi68);
and gate_970(n1061,n393,n1060);
not gate_971(n1062,n1061);
and gate_972(n1063,pi71,n360);
not gate_973(n1064,n1063);
and gate_974(n1065,pi14,n403);
not gate_975(n1066,n1065);
and gate_976(n1067,n1064,n1066);
not gate_977(n1068,n1067);
and gate_978(n1069,n408,n1068);
not gate_979(n1070,n1069);
and gate_980(n1071,n1062,n1070);
not gate_981(n1072,n1071);
and gate_982(n1073,n470,n1071);
not gate_983(n1074,n1073);
and gate_984(n1075,n471,n1072);
not gate_985(n1076,n1075);
and gate_986(n1077,n1074,n1076);
not gate_987(n1078,n1077);
and gate_988(n1079,n1058,n1078);
not gate_989(n1080,n1079);
and gate_990(n1081,n1059,n1077);
not gate_991(n1082,n1081);
and gate_992(n1083,pi15,n97);
not gate_993(n1084,n1083);
and gate_994(n1085,n331,n1084);
not gate_995(n1086,n1085);
and gate_996(n1087,n96,n1086);
and gate_997(n1088,pi71,n1087);
not gate_998(n1089,n1088);
and gate_999(n1090,pi63,n436);
not gate_1000(n1091,n1090);
and gate_1001(n1092,pi31,n439);
not gate_1002(n1093,n1092);
and gate_1003(n1094,n1091,n1093);
not gate_1004(n1095,n1094);
and gate_1005(n1096,n98,n1095);
not gate_1006(n1097,n1096);
and gate_1007(n1098,n1089,n1097);
not gate_1008(n1099,n1098);
and gate_1009(n1100,n95,n1099);
not gate_1010(n1101,n1100);
and gate_1011(n1102,pi47,pi68);
and gate_1012(n1103,n393,n1102);
not gate_1013(n1104,n1103);
and gate_1014(n1105,pi71,n330);
not gate_1015(n1106,n1105);
and gate_1016(n1107,pi15,n403);
not gate_1017(n1108,n1107);
and gate_1018(n1109,n1106,n1108);
not gate_1019(n1110,n1109);
and gate_1020(n1111,n408,n1110);
not gate_1021(n1112,n1111);
and gate_1022(n1113,n1104,n1112);
not gate_1023(n1114,n1113);
and gate_1024(n1115,n470,n1113);
not gate_1025(n1116,n1115);
and gate_1026(n1117,n471,n1114);
not gate_1027(n1118,n1117);
and gate_1028(n1119,n1116,n1118);
not gate_1029(n1120,n1119);
and gate_1030(n1121,n1100,n1120);
not gate_1031(n1122,n1121);
and gate_1032(n1123,n1082,n1121);
not gate_1033(n1124,n1123);
and gate_1034(n1125,n1080,n1124);
and gate_1035(n1126,n1017,n1037);
not gate_1036(n1127,n1126);
and gate_1037(n1128,n1125,n1127);
not gate_1038(n1129,n1128);
and gate_1039(n1130,n1040,n1129);
not gate_1040(n1131,n1130);
and gate_1041(n1132,n997,n1131);
and gate_1042(n1133,n1101,n1119);
not gate_1043(n1134,n1133);
and gate_1044(n1135,n470,n1134);
not gate_1045(n1136,n1135);
and gate_1046(n1137,n1040,n1082);
and gate_1047(n1138,n1135,n1137);
not gate_1048(n1139,n1138);
and gate_1049(n1140,n1132,n1139);
not gate_1050(n1141,n1140);
and gate_1051(n1142,n926,n944);
not gate_1052(n1143,n1142);
and gate_1053(n1144,n1141,n1143);
not gate_1054(n1145,n1144);
and gate_1055(n1146,n865,n907);
and gate_1056(n1147,n1144,n1146);
not gate_1057(n1148,n1147);
and gate_1058(n1149,n957,n1148);
not gate_1059(n1150,n1149);
and gate_1060(n1151,n749,n767);
not gate_1061(n1152,n1151);
and gate_1062(n1153,n1150,n1152);
not gate_1063(n1154,n1153);
and gate_1064(n1155,n690,n730);
and gate_1065(n1156,n1153,n1155);
not gate_1066(n1157,n1156);
and gate_1067(n1158,n782,n1157);
not gate_1068(n1159,n1158);
and gate_1069(n1160,n585,n605);
not gate_1070(n1161,n1160);
and gate_1071(n1162,n1159,n1161);
not gate_1072(n1163,n1162);
and gate_1073(n1164,n607,n1163);
not gate_1074(n1165,n1164);
and gate_1075(n1166,n567,n1165);
not gate_1076(n1167,n1166);
and gate_1077(n1168,n565,n1167);
not gate_1078(n1169,n1168);
and gate_1079(n1170,n525,n1169);
not gate_1080(n1171,n1170);
and gate_1081(n1172,n523,n1171);
not gate_1082(n1173,n1172);
and gate_1083(n1174,n482,n1173);
not gate_1084(n1175,n1174);
and gate_1085(n1176,n483,n1172);
not gate_1086(n1177,n1176);
and gate_1087(n1178,n1175,n1177);
not gate_1088(n1179,n1178);
and gate_1089(n1180,pi66,n94);
not gate_1090(n1181,n1180);
and gate_1091(n1182,n93,pi67);
not gate_1092(n1183,n1182);
and gate_1093(n1184,n1181,n1183);
not gate_1094(n1185,n1184);
and gate_1095(n1186,n1179,n1185);
not gate_1096(n1187,n1186);
and gate_1097(n1188,n428,n1187);
not gate_1098(n1189,n1188);
and gate_1099(n1190,n425,n1189);
not gate_1100(n1191,n1190);
and gate_1101(n1192,n424,n1191);
not gate_1102(po00,n1192);
and gate_1103(n1194,pi72,n101);
not gate_1104(n1195,n1194);
and gate_1105(n1196,n100,pi74);
not gate_1106(n1197,n1196);
and gate_1107(n1198,n1195,n1197);
and gate_1108(n1199,n99,pi73);
not gate_1109(n1200,n1199);
and gate_1110(n1201,n1198,n1200);
not gate_1111(n1202,n1201);
and gate_1112(n1203,n412,n1202);
not gate_1113(n1204,n1203);
and gate_1114(n1205,pi49,pi68);
and gate_1115(n1206,n393,n1205);
not gate_1116(n1207,n1206);
and gate_1117(n1208,pi49,pi70);
and gate_1118(n1209,pi71,n1208);
not gate_1119(n1210,n1209);
and gate_1120(n1211,pi17,n403);
not gate_1121(n1212,n1211);
and gate_1122(n1213,n1210,n1212);
not gate_1123(n1214,n1213);
and gate_1124(n1215,n408,n1214);
not gate_1125(n1216,n1215);
and gate_1126(n1217,n1207,n1216);
not gate_1127(n1218,n1217);
and gate_1128(n1219,n1201,n1218);
not gate_1129(n1220,n1219);
and gate_1130(n1221,n1204,n1220);
not gate_1131(n1222,n1221);
and gate_1132(n1223,pi65,n1222);
not gate_1133(n1224,n1223);
and gate_1134(n1225,n133,n387);
not gate_1135(n1226,n1225);
and gate_1136(n1227,n389,n1226);
and gate_1137(n1228,n92,n1227);
not gate_1138(n1229,n1228);
and gate_1139(n1230,n1224,n1229);
not gate_1140(n1231,n1230);
and gate_1141(n1232,n103,n1231);
not gate_1142(n1233,n1232);
and gate_1143(n1234,n104,n1227);
not gate_1144(n1235,n1234);
and gate_1145(n1236,n1233,n1235);
not gate_1146(n1237,n1236);
and gate_1147(n1238,n91,n1237);
not gate_1148(n1239,n1238);
and gate_1149(n1240,n102,n1222);
not gate_1150(n1241,n1240);
and gate_1151(n1242,n523,n525);
not gate_1152(n1243,n1242);
and gate_1153(n1244,n1168,n1242);
not gate_1154(n1245,n1244);
and gate_1155(n1246,n1169,n1243);
not gate_1156(n1247,n1246);
and gate_1157(n1248,n1245,n1247);
not gate_1158(n1249,n1248);
and gate_1159(n1250,n1185,n1249);
not gate_1160(n1251,n1250);
and gate_1161(n1252,n1241,n1251);
not gate_1162(n1253,n1252);
and gate_1163(n1254,n425,n1253);
not gate_1164(n1255,n1254);
and gate_1165(n1256,n1239,n1255);
not gate_1166(po01,n1256);
and gate_1167(n1258,pi50,pi68);
and gate_1168(n1259,n393,n1258);
not gate_1169(n1260,n1259);
and gate_1170(n1261,pi50,pi70);
and gate_1171(n1262,pi71,n1261);
not gate_1172(n1263,n1262);
and gate_1173(n1264,pi18,n403);
not gate_1174(n1265,n1264);
and gate_1175(n1266,n1263,n1265);
not gate_1176(n1267,n1266);
and gate_1177(n1268,n408,n1267);
not gate_1178(n1269,n1268);
and gate_1179(n1270,n1260,n1269);
not gate_1180(n1271,n1270);
and gate_1181(n1272,n101,n1271);
not gate_1182(n1273,n1272);
and gate_1183(n1274,pi74,n1218);
not gate_1184(n1275,n1274);
and gate_1185(n1276,n1273,n1275);
not gate_1186(n1277,n1276);
and gate_1187(n1278,n99,n100);
not gate_1188(n1279,n1278);
and gate_1189(n1280,n1277,n1278);
not gate_1190(n1281,n1280);
and gate_1191(n1282,n412,n1279);
and gate_1192(n1283,pi72,pi74);
and gate_1193(n1284,pi73,n1283);
not gate_1194(n1285,n1284);
and gate_1195(n1286,n1282,n1285);
not gate_1196(n1287,n1286);
and gate_1197(n1288,n1281,n1287);
and gate_1198(n1289,pi73,n1271);
not gate_1199(n1290,n1289);
and gate_1200(n1291,n1283,n1289);
not gate_1201(n1292,n1291);
and gate_1202(n1293,n1288,n1292);
not gate_1203(n1294,n1293);
and gate_1204(n1295,pi65,n1294);
not gate_1205(n1296,n1295);
and gate_1206(n1297,n150,n385);
not gate_1207(n1298,n1297);
and gate_1208(n1299,n387,n1298);
and gate_1209(n1300,n92,n1299);
not gate_1210(n1301,n1300);
and gate_1211(n1302,n1296,n1301);
not gate_1212(n1303,n1302);
and gate_1213(n1304,n103,n1303);
not gate_1214(n1305,n1304);
and gate_1215(n1306,n104,n1299);
not gate_1216(n1307,n1306);
and gate_1217(n1308,n1305,n1307);
not gate_1218(n1309,n1308);
and gate_1219(n1310,n91,n1309);
not gate_1220(n1311,n1310);
and gate_1221(n1312,n102,n1294);
not gate_1222(n1313,n1312);
and gate_1223(n1314,n565,n567);
not gate_1224(n1315,n1314);
and gate_1225(n1316,n1164,n1314);
not gate_1226(n1317,n1316);
and gate_1227(n1318,n1165,n1315);
not gate_1228(n1319,n1318);
and gate_1229(n1320,n1317,n1319);
not gate_1230(n1321,n1320);
and gate_1231(n1322,n1185,n1321);
not gate_1232(n1323,n1322);
and gate_1233(n1324,n1313,n1323);
not gate_1234(n1325,n1324);
and gate_1235(n1326,n425,n1325);
not gate_1236(n1327,n1326);
and gate_1237(n1328,n1311,n1327);
not gate_1238(po02,n1328);
and gate_1239(n1330,pi51,pi68);
and gate_1240(n1331,n393,n1330);
not gate_1241(n1332,n1331);
and gate_1242(n1333,pi51,pi70);
and gate_1243(n1334,pi71,n1333);
not gate_1244(n1335,n1334);
and gate_1245(n1336,pi19,n403);
not gate_1246(n1337,n1336);
and gate_1247(n1338,n1335,n1337);
not gate_1248(n1339,n1338);
and gate_1249(n1340,n408,n1339);
not gate_1250(n1341,n1340);
and gate_1251(n1342,n1332,n1341);
not gate_1252(n1343,n1342);
and gate_1253(n1344,pi73,pi74);
not gate_1254(n1345,n1344);
and gate_1255(n1346,n1343,n1344);
not gate_1256(n1347,n1346);
and gate_1257(n1348,n412,n1345);
not gate_1258(n1349,n1348);
and gate_1259(n1350,n1347,n1349);
not gate_1260(n1351,n1350);
and gate_1261(n1352,pi72,n1351);
not gate_1262(n1353,n1352);
and gate_1263(n1354,n1196,n1271);
not gate_1264(n1355,n1354);
and gate_1265(n1356,n412,n1344);
not gate_1266(n1357,n1356);
and gate_1267(n1358,n1355,n1357);
and gate_1268(n1359,n100,n1343);
not gate_1269(n1360,n1359);
and gate_1270(n1361,pi73,n1218);
not gate_1271(n1362,n1361);
and gate_1272(n1363,n1360,n1362);
not gate_1273(n1364,n1363);
and gate_1274(n1365,n101,n1364);
not gate_1275(n1366,n1365);
and gate_1276(n1367,n1358,n1366);
not gate_1277(n1368,n1367);
and gate_1278(n1369,n99,n1368);
not gate_1279(n1370,n1369);
and gate_1280(n1371,n1353,n1370);
not gate_1281(n1372,n1371);
and gate_1282(n1373,n102,n1372);
not gate_1283(n1374,n1373);
and gate_1284(n1375,n607,n1161);
not gate_1285(n1376,n1375);
and gate_1286(n1377,n1158,n1375);
not gate_1287(n1378,n1377);
and gate_1288(n1379,n1159,n1376);
not gate_1289(n1380,n1379);
and gate_1290(n1381,n1378,n1380);
not gate_1291(n1382,n1381);
and gate_1292(n1383,n1185,n1382);
not gate_1293(n1384,n1383);
and gate_1294(n1385,n1374,n1384);
not gate_1295(n1386,n1385);
and gate_1296(n1387,n425,n1386);
not gate_1297(n1388,n1387);
and gate_1298(n1389,pi65,n1372);
not gate_1299(n1390,n1389);
and gate_1300(n1391,n168,n383);
not gate_1301(n1392,n1391);
and gate_1302(n1393,n167,n382);
not gate_1303(n1394,n1393);
and gate_1304(n1395,n1392,n1394);
not gate_1305(n1396,n1395);
and gate_1306(n1397,n92,n1396);
not gate_1307(n1398,n1397);
and gate_1308(n1399,n1390,n1398);
not gate_1309(n1400,n1399);
and gate_1310(n1401,n103,n1400);
not gate_1311(n1402,n1401);
and gate_1312(n1403,n104,n1396);
not gate_1313(n1404,n1403);
and gate_1314(n1405,n1402,n1404);
not gate_1315(n1406,n1405);
and gate_1316(n1407,n91,n1406);
not gate_1317(n1408,n1407);
and gate_1318(n1409,n1388,n1408);
not gate_1319(po03,n1409);
and gate_1320(n1411,pi72,n412);
not gate_1321(n1412,n1411);
and gate_1322(n1413,n1345,n1411);
not gate_1323(n1414,n1413);
and gate_1324(n1415,n1196,n1343);
not gate_1325(n1416,n1415);
and gate_1326(n1417,pi52,pi68);
and gate_1327(n1418,n393,n1417);
not gate_1328(n1419,n1418);
and gate_1329(n1420,pi52,pi70);
and gate_1330(n1421,pi71,n1420);
not gate_1331(n1422,n1421);
and gate_1332(n1423,pi20,n403);
not gate_1333(n1424,n1423);
and gate_1334(n1425,n1422,n1424);
not gate_1335(n1426,n1425);
and gate_1336(n1427,n408,n1426);
not gate_1337(n1428,n1427);
and gate_1338(n1429,n1419,n1428);
not gate_1339(n1430,n1429);
and gate_1340(n1431,n100,n1430);
not gate_1341(n1432,n1431);
and gate_1342(n1433,n1290,n1432);
not gate_1343(n1434,n1433);
and gate_1344(n1435,n101,n1434);
not gate_1345(n1436,n1435);
and gate_1346(n1437,n1416,n1436);
not gate_1347(n1438,n1437);
and gate_1348(n1439,n99,n1438);
not gate_1349(n1440,n1439);
and gate_1350(n1441,n1414,n1440);
and gate_1351(n1442,n99,n1218);
not gate_1352(n1443,n1442);
and gate_1353(n1444,pi72,n1430);
not gate_1354(n1445,n1444);
and gate_1355(n1446,n1443,n1445);
not gate_1356(n1447,n1446);
and gate_1357(n1448,n1344,n1447);
not gate_1358(n1449,n1448);
and gate_1359(n1450,n1441,n1449);
not gate_1360(n1451,n1450);
and gate_1361(n1452,pi65,n1451);
not gate_1362(n1453,n1452);
and gate_1363(n1454,n291,n381);
not gate_1364(n1455,n1454);
and gate_1365(n1456,n290,n380);
not gate_1366(n1457,n1456);
and gate_1367(n1458,n1455,n1457);
not gate_1368(n1459,n1458);
and gate_1369(n1460,n92,n1459);
not gate_1370(n1461,n1460);
and gate_1371(n1462,n1453,n1461);
not gate_1372(n1463,n1462);
and gate_1373(n1464,n103,n1463);
not gate_1374(n1465,n1464);
and gate_1375(n1466,n104,n1459);
not gate_1376(n1467,n1466);
and gate_1377(n1468,n1465,n1467);
not gate_1378(n1469,n1468);
and gate_1379(n1470,n91,n1469);
not gate_1380(n1471,n1470);
and gate_1381(n1472,n102,n1451);
not gate_1382(n1473,n1472);
and gate_1383(n1474,n770,n1154);
not gate_1384(n1475,n1474);
and gate_1385(n1476,n730,n1475);
not gate_1386(n1477,n1476);
and gate_1387(n1478,n774,n1477);
not gate_1388(n1479,n1478);
and gate_1389(n1480,n689,n1479);
not gate_1390(n1481,n1480);
and gate_1391(n1482,n777,n1481);
not gate_1392(n1483,n1482);
and gate_1393(n1484,n647,n649);
not gate_1394(n1485,n1484);
and gate_1395(n1486,n1482,n1484);
not gate_1396(n1487,n1486);
and gate_1397(n1488,n1483,n1485);
not gate_1398(n1489,n1488);
and gate_1399(n1490,n1487,n1489);
not gate_1400(n1491,n1490);
and gate_1401(n1492,n1185,n1491);
not gate_1402(n1493,n1492);
and gate_1403(n1494,n1473,n1493);
not gate_1404(n1495,n1494);
and gate_1405(n1496,n425,n1495);
not gate_1406(n1497,n1496);
and gate_1407(n1498,n1471,n1497);
not gate_1408(po04,n1498);
and gate_1409(n1500,pi53,pi68);
and gate_1410(n1501,n393,n1500);
not gate_1411(n1502,n1501);
and gate_1412(n1503,pi53,pi70);
and gate_1413(n1504,pi71,n1503);
not gate_1414(n1505,n1504);
and gate_1415(n1506,pi21,n403);
not gate_1416(n1507,n1506);
and gate_1417(n1508,n1505,n1507);
not gate_1418(n1509,n1508);
and gate_1419(n1510,n408,n1509);
not gate_1420(n1511,n1510);
and gate_1421(n1512,n1502,n1511);
not gate_1422(n1513,n1512);
and gate_1423(n1514,pi72,n1513);
not gate_1424(n1515,n1514);
and gate_1425(n1516,n99,n1271);
not gate_1426(n1517,n1516);
and gate_1427(n1518,n1515,n1517);
not gate_1428(n1519,n1518);
and gate_1429(n1520,pi73,n1519);
not gate_1430(n1521,n1520);
and gate_1431(n1522,n99,n1430);
not gate_1432(n1523,n1522);
and gate_1433(n1524,n1412,n1523);
not gate_1434(n1525,n1524);
and gate_1435(n1526,n100,n1525);
not gate_1436(n1527,n1526);
and gate_1437(n1528,n1521,n1527);
not gate_1438(n1529,n1528);
and gate_1439(n1530,pi74,n1529);
not gate_1440(n1531,n1530);
and gate_1441(n1532,n99,n1343);
not gate_1442(n1533,n1532);
and gate_1443(n1534,n1412,n1533);
not gate_1444(n1535,n1534);
and gate_1445(n1536,pi73,n1535);
not gate_1446(n1537,n1536);
and gate_1447(n1538,n99,n1513);
not gate_1448(n1539,n1538);
and gate_1449(n1540,pi72,n1218);
not gate_1450(n1541,n1540);
and gate_1451(n1542,n1539,n1541);
not gate_1452(n1543,n1542);
and gate_1453(n1544,n100,n1543);
not gate_1454(n1545,n1544);
and gate_1455(n1546,n1537,n1545);
not gate_1456(n1547,n1546);
and gate_1457(n1548,n101,n1547);
not gate_1458(n1549,n1548);
and gate_1459(n1550,n1531,n1549);
not gate_1460(n1551,n1550);
and gate_1461(n1552,pi65,n1551);
not gate_1462(n1553,n1552);
and gate_1463(n1554,n256,n381);
not gate_1464(n1555,n1554);
and gate_1465(n1556,n255,n380);
not gate_1466(n1557,n1556);
and gate_1467(n1558,n1555,n1557);
not gate_1468(n1559,n1558);
and gate_1469(n1560,n92,n1559);
not gate_1470(n1561,n1560);
and gate_1471(n1562,n1553,n1561);
not gate_1472(n1563,n1562);
and gate_1473(n1564,n103,n1563);
not gate_1474(n1565,n1564);
and gate_1475(n1566,n104,n1559);
not gate_1476(n1567,n1566);
and gate_1477(n1568,n1565,n1567);
not gate_1478(n1569,n1568);
and gate_1479(n1570,n91,n1569);
not gate_1480(n1571,n1570);
and gate_1481(n1572,n102,n1551);
not gate_1482(n1573,n1572);
and gate_1483(n1574,n689,n777);
not gate_1484(n1575,n1574);
and gate_1485(n1576,n1478,n1574);
not gate_1486(n1577,n1576);
and gate_1487(n1578,n1479,n1575);
not gate_1488(n1579,n1578);
and gate_1489(n1580,n1577,n1579);
not gate_1490(n1581,n1580);
and gate_1491(n1582,n1185,n1581);
not gate_1492(n1583,n1582);
and gate_1493(n1584,n1573,n1583);
not gate_1494(n1585,n1584);
and gate_1495(n1586,n425,n1585);
not gate_1496(n1587,n1586);
and gate_1497(n1588,n1571,n1587);
not gate_1498(po05,n1588);
and gate_1499(n1590,pi54,pi68);
and gate_1500(n1591,n393,n1590);
not gate_1501(n1592,n1591);
and gate_1502(n1593,pi54,pi70);
and gate_1503(n1594,pi71,n1593);
not gate_1504(n1595,n1594);
and gate_1505(n1596,pi22,n403);
not gate_1506(n1597,n1596);
and gate_1507(n1598,n1595,n1597);
not gate_1508(n1599,n1598);
and gate_1509(n1600,n408,n1599);
not gate_1510(n1601,n1600);
and gate_1511(n1602,n1592,n1601);
not gate_1512(n1603,n1602);
and gate_1513(n1604,pi72,n1603);
not gate_1514(n1605,n1604);
and gate_1515(n1606,n1533,n1605);
not gate_1516(n1607,n1606);
and gate_1517(n1608,pi73,n1607);
not gate_1518(n1609,n1608);
and gate_1519(n1610,n1545,n1609);
not gate_1520(n1611,n1610);
and gate_1521(n1612,pi74,n1611);
not gate_1522(n1613,n1612);
and gate_1523(n1614,pi73,n1525);
not gate_1524(n1615,n1614);
and gate_1525(n1616,n99,n1603);
not gate_1526(n1617,n1616);
and gate_1527(n1618,pi72,n1271);
not gate_1528(n1619,n1618);
and gate_1529(n1620,n1617,n1619);
not gate_1530(n1621,n1620);
and gate_1531(n1622,n100,n1621);
not gate_1532(n1623,n1622);
and gate_1533(n1624,n1615,n1623);
not gate_1534(n1625,n1624);
and gate_1535(n1626,n101,n1625);
not gate_1536(n1627,n1626);
and gate_1537(n1628,n1613,n1627);
not gate_1538(n1629,n1628);
and gate_1539(n1630,pi65,n1629);
not gate_1540(n1631,n1630);
and gate_1541(n1632,n273,n381);
not gate_1542(n1633,n1632);
and gate_1543(n1634,n272,n380);
not gate_1544(n1635,n1634);
and gate_1545(n1636,n1633,n1635);
not gate_1546(n1637,n1636);
and gate_1547(n1638,n92,n1637);
not gate_1548(n1639,n1638);
and gate_1549(n1640,n1631,n1639);
not gate_1550(n1641,n1640);
and gate_1551(n1642,n103,n1641);
not gate_1552(n1643,n1642);
and gate_1553(n1644,n104,n1637);
not gate_1554(n1645,n1644);
and gate_1555(n1646,n1643,n1645);
not gate_1556(n1647,n1646);
and gate_1557(n1648,n91,n1647);
not gate_1558(n1649,n1648);
and gate_1559(n1650,n102,n1629);
not gate_1560(n1651,n1650);
and gate_1561(n1652,n730,n774);
not gate_1562(n1653,n1652);
and gate_1563(n1654,n1474,n1652);
not gate_1564(n1655,n1654);
and gate_1565(n1656,n1475,n1653);
not gate_1566(n1657,n1656);
and gate_1567(n1658,n1655,n1657);
not gate_1568(n1659,n1658);
and gate_1569(n1660,n1185,n1659);
not gate_1570(n1661,n1660);
and gate_1571(n1662,n1651,n1661);
not gate_1572(n1663,n1662);
and gate_1573(n1664,n425,n1663);
not gate_1574(n1665,n1664);
and gate_1575(n1666,n1649,n1665);
not gate_1576(po06,n1666);
and gate_1577(n1668,pi55,pi68);
and gate_1578(n1669,n393,n1668);
not gate_1579(n1670,n1669);
and gate_1580(n1671,pi55,pi70);
and gate_1581(n1672,pi71,n1671);
not gate_1582(n1673,n1672);
and gate_1583(n1674,pi23,n403);
not gate_1584(n1675,n1674);
and gate_1585(n1676,n1673,n1675);
not gate_1586(n1677,n1676);
and gate_1587(n1678,n408,n1677);
not gate_1588(n1679,n1678);
and gate_1589(n1680,n1670,n1679);
not gate_1590(n1681,n1680);
and gate_1591(n1682,pi72,n1681);
not gate_1592(n1683,n1682);
and gate_1593(n1684,n1523,n1683);
not gate_1594(n1685,n1684);
and gate_1595(n1686,pi73,n1685);
not gate_1596(n1687,n1686);
and gate_1597(n1688,n1623,n1687);
not gate_1598(n1689,n1688);
and gate_1599(n1690,pi74,n1689);
not gate_1600(n1691,n1690);
and gate_1601(n1692,n1412,n1539);
not gate_1602(n1693,n1692);
and gate_1603(n1694,pi73,n1693);
not gate_1604(n1695,n1694);
and gate_1605(n1696,n99,n1681);
not gate_1606(n1697,n1696);
and gate_1607(n1698,pi72,n1343);
not gate_1608(n1699,n1698);
and gate_1609(n1700,n1697,n1699);
not gate_1610(n1701,n1700);
and gate_1611(n1702,n100,n1701);
not gate_1612(n1703,n1702);
and gate_1613(n1704,n1695,n1703);
not gate_1614(n1705,n1704);
and gate_1615(n1706,n101,n1705);
not gate_1616(n1707,n1706);
and gate_1617(n1708,n1691,n1707);
not gate_1618(n1709,n1708);
and gate_1619(n1710,n102,n1709);
not gate_1620(n1711,n1710);
and gate_1621(n1712,n770,n1152);
not gate_1622(n1713,n1712);
and gate_1623(n1714,n1149,n1712);
not gate_1624(n1715,n1714);
and gate_1625(n1716,n1150,n1713);
not gate_1626(n1717,n1716);
and gate_1627(n1718,n1715,n1717);
not gate_1628(n1719,n1718);
and gate_1629(n1720,n1185,n1719);
not gate_1630(n1721,n1720);
and gate_1631(n1722,n1711,n1721);
not gate_1632(n1723,n1722);
and gate_1633(n1724,n425,n1723);
not gate_1634(n1725,n1724);
and gate_1635(n1726,pi65,n1709);
not gate_1636(n1727,n1726);
and gate_1637(n1728,n308,n381);
not gate_1638(n1729,n1728);
and gate_1639(n1730,n307,n380);
not gate_1640(n1731,n1730);
and gate_1641(n1732,n1729,n1731);
not gate_1642(n1733,n1732);
and gate_1643(n1734,n92,n1733);
not gate_1644(n1735,n1734);
and gate_1645(n1736,n1727,n1735);
not gate_1646(n1737,n1736);
and gate_1647(n1738,n103,n1737);
not gate_1648(n1739,n1738);
and gate_1649(n1740,n104,n1733);
not gate_1650(n1741,n1740);
and gate_1651(n1742,n1739,n1741);
not gate_1652(n1743,n1742);
and gate_1653(n1744,n91,n1743);
not gate_1654(n1745,n1744);
and gate_1655(n1746,n1725,n1745);
not gate_1656(po07,n1746);
and gate_1657(n1748,pi56,pi68);
and gate_1658(n1749,n393,n1748);
not gate_1659(n1750,n1749);
and gate_1660(n1751,pi56,pi70);
and gate_1661(n1752,pi71,n1751);
not gate_1662(n1753,n1752);
and gate_1663(n1754,pi24,n403);
not gate_1664(n1755,n1754);
and gate_1665(n1756,n1753,n1755);
not gate_1666(n1757,n1756);
and gate_1667(n1758,n408,n1757);
not gate_1668(n1759,n1758);
and gate_1669(n1760,n1750,n1759);
not gate_1670(n1761,n1760);
and gate_1671(n1762,pi72,n1761);
not gate_1672(n1763,n1762);
and gate_1673(n1764,n1539,n1763);
not gate_1674(n1765,n1764);
and gate_1675(n1766,pi73,n1765);
not gate_1676(n1767,n1766);
and gate_1677(n1768,n1703,n1767);
not gate_1678(n1769,n1768);
and gate_1679(n1770,pi74,n1769);
not gate_1680(n1771,n1770);
and gate_1681(n1772,n1412,n1617);
not gate_1682(n1773,n1772);
and gate_1683(n1774,pi73,n1773);
not gate_1684(n1775,n1774);
and gate_1685(n1776,n99,n1761);
not gate_1686(n1777,n1776);
and gate_1687(n1778,n1445,n1777);
not gate_1688(n1779,n1778);
and gate_1689(n1780,n100,n1779);
not gate_1690(n1781,n1780);
and gate_1691(n1782,n1775,n1781);
not gate_1692(n1783,n1782);
and gate_1693(n1784,n101,n1783);
not gate_1694(n1785,n1784);
and gate_1695(n1786,n1771,n1785);
not gate_1696(n1787,n1786);
and gate_1697(n1788,pi65,n1787);
not gate_1698(n1789,n1788);
and gate_1699(n1790,n237,n378);
not gate_1700(n1791,n1790);
and gate_1701(n1792,n203,n1790);
not gate_1702(n1793,n1792);
and gate_1703(n1794,n220,n1793);
not gate_1704(n1795,n1794);
and gate_1705(n1796,n219,n1792);
not gate_1706(n1797,n1796);
and gate_1707(n1798,n1795,n1797);
not gate_1708(n1799,n1798);
and gate_1709(n1800,n92,n1799);
not gate_1710(n1801,n1800);
and gate_1711(n1802,n1789,n1801);
not gate_1712(n1803,n1802);
and gate_1713(n1804,n103,n1803);
not gate_1714(n1805,n1804);
and gate_1715(n1806,n104,n1799);
not gate_1716(n1807,n1806);
and gate_1717(n1808,n1805,n1807);
not gate_1718(n1809,n1808);
and gate_1719(n1810,n91,n1809);
not gate_1720(n1811,n1810);
and gate_1721(n1812,n102,n1787);
not gate_1722(n1813,n1812);
and gate_1723(n1814,n947,n1145);
not gate_1724(n1815,n1814);
and gate_1725(n1816,n907,n1815);
not gate_1726(n1817,n1816);
and gate_1727(n1818,n905,n1817);
not gate_1728(n1819,n1818);
and gate_1729(n1820,n864,n1819);
not gate_1730(n1821,n1820);
and gate_1731(n1822,n952,n1821);
not gate_1732(n1823,n1822);
and gate_1733(n1824,n822,n824);
not gate_1734(n1825,n1824);
and gate_1735(n1826,n1822,n1824);
not gate_1736(n1827,n1826);
and gate_1737(n1828,n1823,n1825);
not gate_1738(n1829,n1828);
and gate_1739(n1830,n1827,n1829);
not gate_1740(n1831,n1830);
and gate_1741(n1832,n1185,n1831);
not gate_1742(n1833,n1832);
and gate_1743(n1834,n1813,n1833);
not gate_1744(n1835,n1834);
and gate_1745(n1836,n425,n1835);
not gate_1746(n1837,n1836);
and gate_1747(n1838,n1811,n1837);
not gate_1748(po08,n1838);
and gate_1749(n1840,pi57,pi68);
and gate_1750(n1841,n393,n1840);
not gate_1751(n1842,n1841);
and gate_1752(n1843,pi57,pi70);
and gate_1753(n1844,pi71,n1843);
not gate_1754(n1845,n1844);
and gate_1755(n1846,pi25,n403);
not gate_1756(n1847,n1846);
and gate_1757(n1848,n1845,n1847);
not gate_1758(n1849,n1848);
and gate_1759(n1850,n408,n1849);
not gate_1760(n1851,n1850);
and gate_1761(n1852,n1842,n1851);
not gate_1762(n1853,n1852);
and gate_1763(n1854,pi72,n1853);
not gate_1764(n1855,n1854);
and gate_1765(n1856,n1617,n1855);
not gate_1766(n1857,n1856);
and gate_1767(n1858,pi73,n1857);
not gate_1768(n1859,n1858);
and gate_1769(n1860,n1781,n1859);
not gate_1770(n1861,n1860);
and gate_1771(n1862,pi74,n1861);
not gate_1772(n1863,n1862);
and gate_1773(n1864,n1541,n1697);
not gate_1774(n1865,n1864);
and gate_1775(n1866,pi73,n1865);
not gate_1776(n1867,n1866);
and gate_1777(n1868,n99,n1853);
not gate_1778(n1869,n1868);
and gate_1779(n1870,n1515,n1869);
not gate_1780(n1871,n1870);
and gate_1781(n1872,n100,n1871);
not gate_1782(n1873,n1872);
and gate_1783(n1874,n1867,n1873);
not gate_1784(n1875,n1874);
and gate_1785(n1876,n101,n1875);
not gate_1786(n1877,n1876);
and gate_1787(n1878,n1863,n1877);
not gate_1788(n1879,n1878);
and gate_1789(n1880,pi65,n1879);
not gate_1790(n1881,n1880);
and gate_1791(n1882,n202,n1790);
not gate_1792(n1883,n1882);
and gate_1793(n1884,n185,n1883);
not gate_1794(n1885,n1884);
and gate_1795(n1886,n184,n1882);
not gate_1796(n1887,n1886);
and gate_1797(n1888,n1885,n1887);
not gate_1798(n1889,n1888);
and gate_1799(n1890,n92,n1889);
not gate_1800(n1891,n1890);
and gate_1801(n1892,n1881,n1891);
not gate_1802(n1893,n1892);
and gate_1803(n1894,n103,n1893);
not gate_1804(n1895,n1894);
and gate_1805(n1896,n104,n1889);
not gate_1806(n1897,n1896);
and gate_1807(n1898,n1895,n1897);
not gate_1808(n1899,n1898);
and gate_1809(n1900,n91,n1899);
not gate_1810(n1901,n1900);
and gate_1811(n1902,n102,n1879);
not gate_1812(n1903,n1902);
and gate_1813(n1904,n864,n952);
not gate_1814(n1905,n1904);
and gate_1815(n1906,n1818,n1904);
not gate_1816(n1907,n1906);
and gate_1817(n1908,n1819,n1905);
not gate_1818(n1909,n1908);
and gate_1819(n1910,n1907,n1909);
not gate_1820(n1911,n1910);
and gate_1821(n1912,n1185,n1911);
not gate_1822(n1913,n1912);
and gate_1823(n1914,n1903,n1913);
not gate_1824(n1915,n1914);
and gate_1825(n1916,n425,n1915);
not gate_1826(n1917,n1916);
and gate_1827(n1918,n1901,n1917);
not gate_1828(po09,n1918);
and gate_1829(n1920,pi58,pi68);
and gate_1830(n1921,n393,n1920);
not gate_1831(n1922,n1921);
and gate_1832(n1923,pi58,pi70);
and gate_1833(n1924,pi71,n1923);
not gate_1834(n1925,n1924);
and gate_1835(n1926,pi26,n403);
not gate_1836(n1927,n1926);
and gate_1837(n1928,n1925,n1927);
not gate_1838(n1929,n1928);
and gate_1839(n1930,n408,n1929);
not gate_1840(n1931,n1930);
and gate_1841(n1932,n1922,n1931);
not gate_1842(n1933,n1932);
and gate_1843(n1934,pi72,n1933);
not gate_1844(n1935,n1934);
and gate_1845(n1936,n1697,n1935);
not gate_1846(n1937,n1936);
and gate_1847(n1938,pi73,n1937);
not gate_1848(n1939,n1938);
and gate_1849(n1940,n1873,n1939);
not gate_1850(n1941,n1940);
and gate_1851(n1942,pi74,n1941);
not gate_1852(n1943,n1942);
and gate_1853(n1944,n1619,n1777);
not gate_1854(n1945,n1944);
and gate_1855(n1946,pi73,n1945);
not gate_1856(n1947,n1946);
and gate_1857(n1948,n99,n1933);
not gate_1858(n1949,n1948);
and gate_1859(n1950,n1605,n1949);
not gate_1860(n1951,n1950);
and gate_1861(n1952,n100,n1951);
not gate_1862(n1953,n1952);
and gate_1863(n1954,n1947,n1953);
not gate_1864(n1955,n1954);
and gate_1865(n1956,n101,n1955);
not gate_1866(n1957,n1956);
and gate_1867(n1958,n1943,n1957);
not gate_1868(n1959,n1958);
and gate_1869(n1960,pi65,n1959);
not gate_1870(n1961,n1960);
and gate_1871(n1962,n201,n1791);
not gate_1872(n1963,n1962);
and gate_1873(n1964,n1883,n1963);
and gate_1874(n1965,n92,n1964);
not gate_1875(n1966,n1965);
and gate_1876(n1967,n1961,n1966);
not gate_1877(n1968,n1967);
and gate_1878(n1969,n103,n1968);
not gate_1879(n1970,n1969);
and gate_1880(n1971,n104,n1964);
not gate_1881(n1972,n1971);
and gate_1882(n1973,n1970,n1972);
not gate_1883(n1974,n1973);
and gate_1884(n1975,n91,n1974);
not gate_1885(n1976,n1975);
and gate_1886(n1977,n102,n1959);
not gate_1887(n1978,n1977);
and gate_1888(n1979,n905,n907);
not gate_1889(n1980,n1979);
and gate_1890(n1981,n1814,n1979);
not gate_1891(n1982,n1981);
and gate_1892(n1983,n1815,n1980);
not gate_1893(n1984,n1983);
and gate_1894(n1985,n1982,n1984);
not gate_1895(n1986,n1985);
and gate_1896(n1987,n1185,n1986);
not gate_1897(n1988,n1987);
and gate_1898(n1989,n1978,n1988);
not gate_1899(n1990,n1989);
and gate_1900(n1991,n425,n1990);
not gate_1901(n1992,n1991);
and gate_1902(n1993,n1976,n1992);
not gate_1903(po10,n1993);
and gate_1904(n1995,pi59,pi68);
and gate_1905(n1996,n393,n1995);
not gate_1906(n1997,n1996);
and gate_1907(n1998,pi59,pi70);
and gate_1908(n1999,pi71,n1998);
not gate_1909(n2000,n1999);
and gate_1910(n2001,pi27,n403);
not gate_1911(n2002,n2001);
and gate_1912(n2003,n2000,n2002);
not gate_1913(n2004,n2003);
and gate_1914(n2005,n408,n2004);
not gate_1915(n2006,n2005);
and gate_1916(n2007,n1997,n2006);
not gate_1917(n2008,n2007);
and gate_1918(n2009,pi72,n2008);
not gate_1919(n2010,n2009);
and gate_1920(n2011,n1777,n2010);
not gate_1921(n2012,n2011);
and gate_1922(n2013,pi73,n2012);
not gate_1923(n2014,n2013);
and gate_1924(n2015,n1953,n2014);
not gate_1925(n2016,n2015);
and gate_1926(n2017,pi74,n2016);
not gate_1927(n2018,n2017);
and gate_1928(n2019,n1699,n1869);
not gate_1929(n2020,n2019);
and gate_1930(n2021,pi73,n2020);
not gate_1931(n2022,n2021);
and gate_1932(n2023,n99,n2008);
not gate_1933(n2024,n2023);
and gate_1934(n2025,n1683,n2024);
not gate_1935(n2026,n2025);
and gate_1936(n2027,n100,n2026);
not gate_1937(n2028,n2027);
and gate_1938(n2029,n2022,n2028);
not gate_1939(n2030,n2029);
and gate_1940(n2031,n101,n2030);
not gate_1941(n2032,n2031);
and gate_1942(n2033,n2018,n2032);
not gate_1943(n2034,n2033);
and gate_1944(n2035,n102,n2034);
not gate_1945(n2036,n2035);
and gate_1946(n2037,n947,n1143);
not gate_1947(n2038,n2037);
and gate_1948(n2039,n1140,n2037);
not gate_1949(n2040,n2039);
and gate_1950(n2041,n1141,n2038);
not gate_1951(n2042,n2041);
and gate_1952(n2043,n2040,n2042);
not gate_1953(n2044,n2043);
and gate_1954(n2045,n1185,n2044);
not gate_1955(n2046,n2045);
and gate_1956(n2047,n2036,n2046);
not gate_1957(n2048,n2047);
and gate_1958(n2049,n425,n2048);
not gate_1959(n2050,n2049);
and gate_1960(n2051,pi65,n2034);
not gate_1961(n2052,n2051);
and gate_1962(n2053,n236,n379);
not gate_1963(n2054,n2053);
and gate_1964(n2055,n1791,n2054);
and gate_1965(n2056,n92,n2055);
not gate_1966(n2057,n2056);
and gate_1967(n2058,n2052,n2057);
not gate_1968(n2059,n2058);
and gate_1969(n2060,n103,n2059);
not gate_1970(n2061,n2060);
and gate_1971(n2062,n104,n2055);
not gate_1972(n2063,n2062);
and gate_1973(n2064,n2061,n2063);
not gate_1974(n2065,n2064);
and gate_1975(n2066,n91,n2065);
not gate_1976(n2067,n2066);
and gate_1977(n2068,n2050,n2067);
not gate_1978(po11,n2068);
and gate_1979(n2070,pi60,pi68);
and gate_1980(n2071,n393,n2070);
not gate_1981(n2072,n2071);
and gate_1982(n2073,pi60,pi70);
and gate_1983(n2074,pi71,n2073);
not gate_1984(n2075,n2074);
and gate_1985(n2076,pi28,n403);
not gate_1986(n2077,n2076);
and gate_1987(n2078,n2075,n2077);
not gate_1988(n2079,n2078);
and gate_1989(n2080,n408,n2079);
not gate_1990(n2081,n2080);
and gate_1991(n2082,n2072,n2081);
not gate_1992(n2083,n2082);
and gate_1993(n2084,pi72,n2083);
not gate_1994(n2085,n2084);
and gate_1995(n2086,n1869,n2085);
not gate_1996(n2087,n2086);
and gate_1997(n2088,pi73,n2087);
not gate_1998(n2089,n2088);
and gate_1999(n2090,n2028,n2089);
not gate_2000(n2091,n2090);
and gate_2001(n2092,pi74,n2091);
not gate_2002(n2093,n2092);
and gate_2003(n2094,n1445,n1949);
not gate_2004(n2095,n2094);
and gate_2005(n2096,pi73,n2095);
not gate_2006(n2097,n2096);
and gate_2007(n2098,n99,n2083);
not gate_2008(n2099,n2098);
and gate_2009(n2100,n1763,n2099);
not gate_2010(n2101,n2100);
and gate_2011(n2102,n100,n2101);
not gate_2012(n2103,n2102);
and gate_2013(n2104,n2097,n2103);
not gate_2014(n2105,n2104);
and gate_2015(n2106,n101,n2105);
not gate_2016(n2107,n2106);
and gate_2017(n2108,n2093,n2107);
not gate_2018(n2109,n2108);
and gate_2019(n2110,pi65,n2109);
not gate_2020(n2111,n2110);
and gate_2021(n2112,n327,n377);
not gate_2022(n2113,n2112);
and gate_2023(n2114,n326,n376);
not gate_2024(n2115,n2114);
and gate_2025(n2116,n2113,n2115);
not gate_2026(n2117,n2116);
and gate_2027(n2118,n92,n2117);
not gate_2028(n2119,n2118);
and gate_2029(n2120,n2111,n2119);
not gate_2030(n2121,n2120);
and gate_2031(n2122,n103,n2121);
not gate_2032(n2123,n2122);
and gate_2033(n2124,n104,n2117);
not gate_2034(n2125,n2124);
and gate_2035(n2126,n2123,n2125);
not gate_2036(n2127,n2126);
and gate_2037(n2128,n91,n2127);
not gate_2038(n2129,n2128);
and gate_2039(n2130,n102,n2109);
not gate_2040(n2131,n2130);
and gate_2041(n2132,n1122,n1136);
not gate_2042(n2133,n2132);
and gate_2043(n2134,n1082,n2133);
not gate_2044(n2135,n2134);
and gate_2045(n2136,n1080,n2135);
not gate_2046(n2137,n2136);
and gate_2047(n2138,n1039,n2137);
not gate_2048(n2139,n2138);
and gate_2049(n2140,n1127,n2139);
not gate_2050(n2141,n2140);
and gate_2051(n2142,n997,n999);
not gate_2052(n2143,n2142);
and gate_2053(n2144,n2140,n2142);
not gate_2054(n2145,n2144);
and gate_2055(n2146,n2141,n2143);
not gate_2056(n2147,n2146);
and gate_2057(n2148,n2145,n2147);
not gate_2058(n2149,n2148);
and gate_2059(n2150,n1185,n2149);
not gate_2060(n2151,n2150);
and gate_2061(n2152,n2131,n2151);
not gate_2062(n2153,n2152);
and gate_2063(n2154,n425,n2153);
not gate_2064(n2155,n2154);
and gate_2065(n2156,n2129,n2155);
not gate_2066(po12,n2156);
and gate_2067(n2158,pi61,pi68);
and gate_2068(n2159,n393,n2158);
not gate_2069(n2160,n2159);
and gate_2070(n2161,pi61,pi70);
and gate_2071(n2162,pi71,n2161);
not gate_2072(n2163,n2162);
and gate_2073(n2164,pi29,n403);
not gate_2074(n2165,n2164);
and gate_2075(n2166,n2163,n2165);
not gate_2076(n2167,n2166);
and gate_2077(n2168,n408,n2167);
not gate_2078(n2169,n2168);
and gate_2079(n2170,n2160,n2169);
not gate_2080(n2171,n2170);
and gate_2081(n2172,pi72,n2171);
not gate_2082(n2173,n2172);
and gate_2083(n2174,n1949,n2173);
not gate_2084(n2175,n2174);
and gate_2085(n2176,pi73,n2175);
not gate_2086(n2177,n2176);
and gate_2087(n2178,n2103,n2177);
not gate_2088(n2179,n2178);
and gate_2089(n2180,pi74,n2179);
not gate_2090(n2181,n2180);
and gate_2091(n2182,n1515,n2024);
not gate_2092(n2183,n2182);
and gate_2093(n2184,pi73,n2183);
not gate_2094(n2185,n2184);
and gate_2095(n2186,n99,n2171);
not gate_2096(n2187,n2186);
and gate_2097(n2188,n1855,n2187);
not gate_2098(n2189,n2188);
and gate_2099(n2190,n100,n2189);
not gate_2100(n2191,n2190);
and gate_2101(n2192,n2185,n2191);
not gate_2102(n2193,n2192);
and gate_2103(n2194,n101,n2193);
not gate_2104(n2195,n2194);
and gate_2105(n2196,n2181,n2195);
not gate_2106(n2197,n2196);
and gate_2107(n2198,pi65,n2197);
not gate_2108(n2199,n2198);
and gate_2109(n2200,n128,n337);
not gate_2110(n2201,n2200);
and gate_2111(n2202,n340,n2201);
not gate_2112(n2203,n2202);
and gate_2113(n2204,n369,n2203);
not gate_2114(n2205,n2204);
and gate_2115(n2206,n357,n2205);
not gate_2116(n2207,n2206);
and gate_2117(n2208,n356,n2204);
not gate_2118(n2209,n2208);
and gate_2119(n2210,n2207,n2209);
not gate_2120(n2211,n2210);
and gate_2121(n2212,n92,n2211);
not gate_2122(n2213,n2212);
and gate_2123(n2214,n2199,n2213);
not gate_2124(n2215,n2214);
and gate_2125(n2216,n103,n2215);
not gate_2126(n2217,n2216);
and gate_2127(n2218,n104,n2211);
not gate_2128(n2219,n2218);
and gate_2129(n2220,n2217,n2219);
not gate_2130(n2221,n2220);
and gate_2131(n2222,n91,n2221);
not gate_2132(n2223,n2222);
and gate_2133(n2224,n102,n2197);
not gate_2134(n2225,n2224);
and gate_2135(n2226,n1039,n1127);
not gate_2136(n2227,n2226);
and gate_2137(n2228,n2136,n2226);
not gate_2138(n2229,n2228);
and gate_2139(n2230,n2137,n2227);
not gate_2140(n2231,n2230);
and gate_2141(n2232,n2229,n2231);
not gate_2142(n2233,n2232);
and gate_2143(n2234,n1185,n2233);
not gate_2144(n2235,n2234);
and gate_2145(n2236,n2225,n2235);
not gate_2146(n2237,n2236);
and gate_2147(n2238,n425,n2237);
not gate_2148(n2239,n2238);
and gate_2149(n2240,n2223,n2239);
not gate_2150(po13,n2240);
and gate_2151(n2242,pi62,pi68);
and gate_2152(n2243,n393,n2242);
not gate_2153(n2244,n2243);
and gate_2154(n2245,pi62,pi70);
and gate_2155(n2246,pi71,n2245);
not gate_2156(n2247,n2246);
and gate_2157(n2248,pi30,n403);
not gate_2158(n2249,n2248);
and gate_2159(n2250,n2247,n2249);
not gate_2160(n2251,n2250);
and gate_2161(n2252,n408,n2251);
not gate_2162(n2253,n2252);
and gate_2163(n2254,n2244,n2253);
not gate_2164(n2255,n2254);
and gate_2165(n2256,pi72,n2255);
not gate_2166(n2257,n2256);
and gate_2167(n2258,n2024,n2257);
not gate_2168(n2259,n2258);
and gate_2169(n2260,pi73,n2259);
not gate_2170(n2261,n2260);
and gate_2171(n2262,n2191,n2261);
not gate_2172(n2263,n2262);
and gate_2173(n2264,pi74,n2263);
not gate_2174(n2265,n2264);
and gate_2175(n2266,n1605,n2099);
not gate_2176(n2267,n2266);
and gate_2177(n2268,pi73,n2267);
not gate_2178(n2269,n2268);
and gate_2179(n2270,n99,n2255);
not gate_2180(n2271,n2270);
and gate_2181(n2272,n1935,n2271);
not gate_2182(n2273,n2272);
and gate_2183(n2274,n100,n2273);
not gate_2184(n2275,n2274);
and gate_2185(n2276,n2269,n2275);
not gate_2186(n2277,n2276);
and gate_2187(n2278,n101,n2277);
not gate_2188(n2279,n2278);
and gate_2189(n2280,n2265,n2279);
not gate_2190(n2281,n2280);
and gate_2191(n2282,pi65,n2281);
not gate_2192(n2283,n2282);
and gate_2193(n2284,n340,n374);
not gate_2194(n2285,n2284);
and gate_2195(n2286,n339,n373);
not gate_2196(n2287,n2286);
and gate_2197(n2288,n2285,n2287);
not gate_2198(n2289,n2288);
and gate_2199(n2290,n92,n2289);
not gate_2200(n2291,n2290);
and gate_2201(n2292,n2283,n2291);
not gate_2202(n2293,n2292);
and gate_2203(n2294,n103,n2293);
not gate_2204(n2295,n2294);
and gate_2205(n2296,n104,n2289);
not gate_2206(n2297,n2296);
and gate_2207(n2298,n2295,n2297);
not gate_2208(n2299,n2298);
and gate_2209(n2300,n91,n2299);
not gate_2210(n2301,n2300);
and gate_2211(n2302,n102,n2281);
not gate_2212(n2303,n2302);
and gate_2213(n2304,n1080,n1082);
not gate_2214(n2305,n2304);
and gate_2215(n2306,n2132,n2304);
not gate_2216(n2307,n2306);
and gate_2217(n2308,n2133,n2305);
not gate_2218(n2309,n2308);
and gate_2219(n2310,n2307,n2309);
not gate_2220(n2311,n2310);
and gate_2221(n2312,n1185,n2311);
not gate_2222(n2313,n2312);
and gate_2223(n2314,n2303,n2313);
not gate_2224(n2315,n2314);
and gate_2225(n2316,n425,n2315);
not gate_2226(n2317,n2316);
and gate_2227(n2318,n2301,n2317);
not gate_2228(po14,n2318);
and gate_2229(n2320,pi63,pi68);
and gate_2230(n2321,n393,n2320);
not gate_2231(n2322,n2321);
and gate_2232(n2323,pi63,pi70);
and gate_2233(n2324,pi71,n2323);
not gate_2234(n2325,n2324);
and gate_2235(n2326,pi31,n403);
not gate_2236(n2327,n2326);
and gate_2237(n2328,n2325,n2327);
not gate_2238(n2329,n2328);
and gate_2239(n2330,n408,n2329);
not gate_2240(n2331,n2330);
and gate_2241(n2332,n2322,n2331);
not gate_2242(n2333,n2332);
and gate_2243(n2334,pi72,n2333);
not gate_2244(n2335,n2334);
and gate_2245(n2336,n2099,n2335);
not gate_2246(n2337,n2336);
and gate_2247(n2338,pi73,n2337);
not gate_2248(n2339,n2338);
and gate_2249(n2340,n2275,n2339);
not gate_2250(n2341,n2340);
and gate_2251(n2342,pi74,n2341);
not gate_2252(n2343,n2342);
and gate_2253(n2344,n1683,n2187);
not gate_2254(n2345,n2344);
and gate_2255(n2346,pi73,n2345);
not gate_2256(n2347,n2346);
and gate_2257(n2348,n99,n2333);
not gate_2258(n2349,n2348);
and gate_2259(n2350,n2010,n2349);
not gate_2260(n2351,n2350);
and gate_2261(n2352,n100,n2351);
not gate_2262(n2353,n2352);
and gate_2263(n2354,n2347,n2353);
not gate_2264(n2355,n2354);
and gate_2265(n2356,n101,n2355);
not gate_2266(n2357,n2356);
and gate_2267(n2358,n2343,n2357);
not gate_2268(n2359,n2358);
and gate_2269(n2360,pi65,n2359);
not gate_2270(n2361,n2360);
and gate_2271(n2362,n92,n337);
not gate_2272(n2363,n2362);
and gate_2273(n2364,n2361,n2363);
not gate_2274(n2365,n2364);
and gate_2275(n2366,n103,n2365);
not gate_2276(n2367,n2366);
and gate_2277(n2368,n104,n337);
not gate_2278(n2369,n2368);
and gate_2279(n2370,n2367,n2369);
not gate_2280(n2371,n2370);
and gate_2281(n2372,n91,n2371);
not gate_2282(n2373,n2372);
and gate_2283(n2374,n102,n2359);
not gate_2284(n2375,n2374);
and gate_2285(n2376,n1101,n1113);
not gate_2286(n2377,n2376);
and gate_2287(n2378,n1100,n1114);
not gate_2288(n2379,n2378);
and gate_2289(n2380,n2377,n2379);
and gate_2290(n2381,n1185,n2380);
not gate_2291(n2382,n2381);
and gate_2292(n2383,n2375,n2382);
not gate_2293(n2384,n2383);
and gate_2294(n2385,n425,n2384);
not gate_2295(n2386,n2385);
and gate_2296(n2387,n2373,n2386);
not gate_2297(po15,n2387);
endmodule
