// Verilog File 
module i9 (pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
pi39,pi40,pi41,pi42,pi43,pi44,pi45,pi46,pi47,pi48,
pi49,pi50,pi51,pi52,pi53,pi54,pi55,pi56,pi57,pi58,
pi59,pi60,pi61,pi62,pi63,pi64,pi65,pi66,pi67,pi68,
pi69,pi70,pi71,pi72,pi73,pi74,pi75,pi76,pi77,pi78,
pi79,pi80,pi81,pi82,pi83,pi84,pi85,pi86,pi87,po00,
po01,po02,po03,po04,po05,po06,po07,po08,po09,po10,
po11,po12,po13,po14,po15,po16,po17,po18,po19,po20,
po21,po22,po23,po24,po25,po26,po27,po28,po29,po30,
po31,po32,po33,po34,po35,po36,po37,po38,po39,po40,
po41,po42,po43,po44,po45,po46,po47,po48,po49,po50,
po51,po52,po53,po54,po55,po56,po57,po58,po59,po60,
po61,po62);

input pi00,pi01,pi02,pi03,pi04,pi05,pi06,pi07,pi08,
pi09,pi10,pi11,pi12,pi13,pi14,pi15,pi16,pi17,pi18,
pi19,pi20,pi21,pi22,pi23,pi24,pi25,pi26,pi27,pi28,
pi29,pi30,pi31,pi32,pi33,pi34,pi35,pi36,pi37,pi38,
pi39,pi40,pi41,pi42,pi43,pi44,pi45,pi46,pi47,pi48,
pi49,pi50,pi51,pi52,pi53,pi54,pi55,pi56,pi57,pi58,
pi59,pi60,pi61,pi62,pi63,pi64,pi65,pi66,pi67,pi68,
pi69,pi70,pi71,pi72,pi73,pi74,pi75,pi76,pi77,pi78,
pi79,pi80,pi81,pi82,pi83,pi84,pi85,pi86,pi87;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18,
po19,po20,po21,po22,po23,po24,po25,po26,po27,po28,
po29,po30,po31,po32,po33,po34,po35,po36,po37,po38,
po39,po40,po41,po42,po43,po44,po45,po46,po47,po48,
po49,po50,po51,po52,po53,po54,po55,po56,po57,po58,
po59,po60,po61,po62;

wire n151,n152,n153,n154,n155,n156,n157,n158,n159,
n160,n161,n162,n163,n164,n165,n166,n167,n168,n169,
n170,n171,n172,n173,n174,n175,n176,n177,n178,n179,
n180,n181,n182,n183,n184,n185,n186,n187,n188,n189,
n190,n191,n192,n193,n194,n195,n196,n197,n198,n199,
n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,
n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,
n220,n221,n222,n223,n224,n225,n226,n227,n228,n229,
n230,n231,n232,n233,n234,n235,n236,n237,n239,n240,
n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,
n251,n252,n253,n254,n255,n257,n258,n259,n260,n261,
n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,
n272,n273,n275,n276,n277,n278,n279,n280,n281,n282,
n283,n284,n285,n286,n287,n288,n289,n290,n291,n293,
n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,
n304,n305,n306,n307,n308,n309,n311,n312,n313,n314,
n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,
n325,n326,n327,n329,n330,n331,n332,n333,n334,n335,
n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,
n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,
n357,n358,n359,n360,n361,n362,n363,n365,n366,n367,
n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,
n378,n379,n380,n381,n383,n384,n385,n386,n387,n388,
n389,n390,n391,n392,n393,n394,n395,n396,n397,n398,
n399,n401,n402,n403,n404,n405,n406,n407,n408,n409,
n410,n411,n412,n413,n414,n415,n416,n417,n419,n420,
n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,
n431,n432,n433,n435,n436,n437,n438,n439,n440,n441,
n442,n443,n444,n445,n446,n447,n448,n449,n451,n452,
n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,
n463,n464,n465,n467,n468,n469,n470,n471,n472,n473,
n474,n475,n476,n477,n478,n479,n480,n481,n483,n484,
n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,
n495,n496,n497,n499,n500,n501,n502,n503,n504,n505,
n506,n507,n508,n509,n510,n511,n512,n513,n515,n516,
n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,
n527,n528,n529,n531,n532,n533,n534,n535,n536,n537,
n538,n539,n540,n541,n542,n543,n544,n545,n547,n548,
n549,n550,n551,n552,n553,n554,n555,n556,n557,n558,
n559,n560,n561,n563,n564,n565,n566,n567,n568,n569,
n570,n571,n572,n573,n574,n575,n576,n577,n579,n580,
n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,
n591,n592,n593,n595,n596,n597,n598,n599,n600,n601,
n602,n603,n604,n605,n606,n607,n608,n609,n611,n612,
n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,
n623,n624,n625,n627,n628,n629,n630,n631,n632,n633,
n634,n635,n636,n637,n638,n639,n641,n642,n643,n644,
n645,n646,n647,n648,n649,n650,n651,n652,n653,n655,
n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,
n666,n667,n669,n670,n671,n672,n673,n674,n675,n676,
n677,n678,n679,n680,n681,n683,n684,n685,n686,n687,
n688,n689,n690,n691,n692,n693,n694,n695,n697,n698,
n699,n700,n701,n702,n703,n704,n705,n706,n707,n708,
n709,n711,n712,n713,n714,n715,n716,n717,n718,n719,
n720,n721,n722,n723,n725,n726,n727,n728,n729,n730,
n731,n732,n733,n734,n735,n736,n737,n738,n739,n741,
n742,n743,n744,n745,n746,n747,n748,n749,n750,n751,
n752,n753,n754,n755,n757,n758,n759,n760,n761,n762,
n763,n764,n765,n766,n767,n768,n769,n770,n771,n773,
n774,n775,n776,n777,n778,n779,n780,n781,n782,n783,
n784,n785,n786,n787,n789,n790,n791,n792,n793,n794,
n795,n796,n797,n798,n799,n800,n801,n802,n803,n804,
n806,n807,n808,n809,n810,n811,n812,n813,n814,n815,
n816,n817,n818,n819,n821,n822,n823,n824,n825,n826,
n827,n828,n829,n830,n831,n832,n833,n834,n836,n837,
n838,n839,n840,n841,n842,n843,n844,n845,n846,n847,
n849,n850,n851,n852,n853,n854,n855,n856,n857,n858,
n859,n860,n862,n863,n864,n865,n866,n867,n868,n869,
n870,n871,n872,n873,n875,n876,n877,n878,n879,n880,
n881,n882,n883,n884,n885,n886,n888,n889,n890,n891,
n892,n893,n894,n895,n896,n897,n898,n899,n901,n902,
n903,n904,n905,n906,n907,n908,n909,n910,n911,n912,
n914,n915,n916,n917,n918,n919,n920,n921,n922,n923,
n924,n925,n927,n928,n929,n930,n931,n932,n933,n934,
n935,n936,n937,n938,n940,n941,n942,n943,n944,n945,
n946,n947,n948,n949,n950,n951,n953,n954,n955,n956,
n957,n958,n959,n960,n961,n962,n963,n964,n965,n966,
n967,n968,n969,n970,n972,n973,n974,n975,n976,n977,
n978,n979,n980,n981,n982,n983,n984,n985,n986,n987,
n988,n989,n991,n992,n993,n994,n995,n996,n997,n998,
n999,n1000,n1001,n1002,n1003,n1004,n1005,n1006,n1007,n1008,
n1010,n1011,n1012,n1013,n1014,n1015,n1016,n1017,n1018,n1019,
n1020,n1021,n1022,n1023,n1024,n1025,n1026,n1027,n1029,n1030,
n1031,n1032,n1033,n1034,n1035,n1036,n1037,n1038,n1039,n1040,
n1041,n1042,n1043,n1044,n1045,n1046,n1048,n1049,n1050,n1051,
n1052,n1053,n1054,n1055,n1056,n1057,n1058,n1059,n1060,n1061,
n1062,n1063,n1065,n1066,n1067,n1068,n1069,n1070,n1071,n1072,
n1073,n1074,n1075,n1076,n1077,n1078,n1079,n1080,n1082,n1083,
n1084,n1085,n1086,n1087,n1088,n1089,n1090,n1091,n1092,n1093,
n1094,n1095,n1097,n1098,n1099,n1100,n1101,n1102,n1103,n1104,
n1105,n1106,n1107,n1108,n1109,n1110,n1112,n1113,n1114,n1115,
n1116,n1117,n1118,n1119,n1120,n1121,n1122,n1124,n1125,n1126,
n1127,n1128,n1129,n1130,n1131,n1132,n1133,n1134,n1136,n1137,
n1138,n1139,n1140,n1141,n1142,n1143,n1144,n1146,n1147,n1148,
n1149,n1150,n1151,n1152,n1153,n1154,n1156,n1157,n1158,n1159,
n1160,n1161,n1162,n1163,n1164,n1166,n1167,n1168,n1169,n1170,
n1171,n1172,n1173,n1174,n1176,n1177,n1178,n1179,n1180,n1181,
n1182,n1183,n1184;
not gate_0(n151,pi00);
not gate_1(n152,pi01);
not gate_2(n153,pi02);
not gate_3(n154,pi03);
not gate_4(n155,pi04);
not gate_5(n156,pi05);
not gate_6(n157,pi06);
and gate_7(n158,n152,pi03);
and gate_8(n159,n153,n158);
not gate_9(n160,n159);
and gate_10(n161,n152,pi07);
and gate_11(n162,n153,n161);
not gate_12(n163,n162);
and gate_13(n164,n153,n157);
and gate_14(n165,n152,n164);
and gate_15(n166,n156,n165);
not gate_16(n167,n166);
and gate_17(n168,n163,n167);
and gate_18(n169,n160,n168);
and gate_19(n170,n154,n155);
and gate_20(n171,pi07,n170);
not gate_21(n172,n171);
and gate_22(n173,pi01,n154);
and gate_23(n174,pi08,n173);
not gate_24(n175,n174);
and gate_25(n176,n156,n170);
not gate_26(n177,n176);
and gate_27(n178,n154,n156);
and gate_28(n179,pi01,n178);
and gate_29(n180,n164,n179);
not gate_30(n181,n180);
and gate_31(n182,n177,n181);
and gate_32(n183,n175,n182);
and gate_33(n184,n172,n183);
and gate_34(n185,n169,n184);
not gate_35(n186,n185);
and gate_36(n187,pi02,n154);
and gate_37(n188,pi01,n187);
and gate_38(n189,n151,n188);
not gate_39(n190,n189);
and gate_40(n191,n152,n178);
and gate_41(n192,pi04,n191);
and gate_42(n193,pi02,n192);
and gate_43(n194,n157,n193);
not gate_44(n195,n194);
and gate_45(n196,n152,n187);
and gate_46(n197,pi08,n196);
not gate_47(n198,n197);
and gate_48(n199,n195,n198);
and gate_49(n200,n190,n199);
and gate_50(n201,n183,n200);
and gate_51(n202,pi00,pi02);
not gate_52(n203,n202);
and gate_53(n204,n154,n203);
not gate_54(n205,n204);
and gate_55(n206,pi01,n205);
not gate_56(n207,n206);
and gate_57(n208,n172,n207);
and gate_58(n209,pi02,pi03);
not gate_59(n210,n209);
and gate_60(n211,n169,n210);
and gate_61(n212,n208,n211);
and gate_62(n213,n201,n212);
not gate_63(n214,n213);
and gate_64(n215,n169,n200);
not gate_65(n216,n215);
and gate_66(n217,n214,n215);
and gate_67(n218,n186,n217);
not gate_68(n219,n218);
and gate_69(n220,pi17,n218);
not gate_70(n221,n220);
and gate_71(n222,pi09,n185);
not gate_72(n223,n222);
and gate_73(n224,n217,n222);
not gate_74(n225,n224);
and gate_75(n226,n214,n225);
and gate_76(n227,n221,n226);
and gate_77(n228,n214,n216);
and gate_78(n229,pi20,n185);
not gate_79(n230,n229);
and gate_80(n231,pi24,n186);
not gate_81(n232,n231);
and gate_82(n233,n230,n232);
not gate_83(n234,n233);
and gate_84(n235,n228,n234);
not gate_85(n236,n235);
and gate_86(n237,n227,n236);
not gate_87(po00,n237);
and gate_88(n239,pi18,n218);
not gate_89(n240,n239);
and gate_90(n241,pi10,n185);
not gate_91(n242,n241);
and gate_92(n243,n217,n241);
not gate_93(n244,n243);
and gate_94(n245,n214,n244);
and gate_95(n246,n240,n245);
and gate_96(n247,pi21,n185);
not gate_97(n248,n247);
and gate_98(n249,pi25,n186);
not gate_99(n250,n249);
and gate_100(n251,n248,n250);
not gate_101(n252,n251);
and gate_102(n253,n228,n252);
not gate_103(n254,n253);
and gate_104(n255,n246,n254);
not gate_105(po01,n255);
and gate_106(n257,pi19,n218);
not gate_107(n258,n257);
and gate_108(n259,pi11,n185);
not gate_109(n260,n259);
and gate_110(n261,n217,n259);
not gate_111(n262,n261);
and gate_112(n263,n214,n262);
and gate_113(n264,n258,n263);
and gate_114(n265,pi22,n185);
not gate_115(n266,n265);
and gate_116(n267,pi26,n186);
not gate_117(n268,n267);
and gate_118(n269,n266,n268);
not gate_119(n270,n269);
and gate_120(n271,n228,n270);
not gate_121(n272,n271);
and gate_122(n273,n264,n272);
not gate_123(po02,n273);
and gate_124(n275,pi20,n218);
not gate_125(n276,n275);
and gate_126(n277,pi12,n185);
not gate_127(n278,n277);
and gate_128(n279,n217,n277);
not gate_129(n280,n279);
and gate_130(n281,n214,n280);
and gate_131(n282,n276,n281);
and gate_132(n283,pi23,n185);
not gate_133(n284,n283);
and gate_134(n285,pi27,n186);
not gate_135(n286,n285);
and gate_136(n287,n284,n286);
not gate_137(n288,n287);
and gate_138(n289,n228,n288);
not gate_139(n290,n289);
and gate_140(n291,n282,n290);
not gate_141(po03,n291);
and gate_142(n293,pi21,n218);
not gate_143(n294,n293);
and gate_144(n295,pi13,n185);
not gate_145(n296,n295);
and gate_146(n297,n217,n295);
not gate_147(n298,n297);
and gate_148(n299,n214,n298);
and gate_149(n300,n294,n299);
and gate_150(n301,pi24,n185);
not gate_151(n302,n301);
and gate_152(n303,pi28,n186);
not gate_153(n304,n303);
and gate_154(n305,n302,n304);
not gate_155(n306,n305);
and gate_156(n307,n228,n306);
not gate_157(n308,n307);
and gate_158(n309,n300,n308);
not gate_159(po04,n309);
and gate_160(n311,pi22,n218);
not gate_161(n312,n311);
and gate_162(n313,pi14,n185);
not gate_163(n314,n313);
and gate_164(n315,n217,n313);
not gate_165(n316,n315);
and gate_166(n317,n214,n316);
and gate_167(n318,n312,n317);
and gate_168(n319,pi25,n185);
not gate_169(n320,n319);
and gate_170(n321,pi29,n186);
not gate_171(n322,n321);
and gate_172(n323,n320,n322);
not gate_173(n324,n323);
and gate_174(n325,n228,n324);
not gate_175(n326,n325);
and gate_176(n327,n318,n326);
not gate_177(po05,n327);
and gate_178(n329,pi23,n218);
not gate_179(n330,n329);
and gate_180(n331,pi15,n185);
not gate_181(n332,n331);
and gate_182(n333,n217,n331);
not gate_183(n334,n333);
and gate_184(n335,n214,n334);
and gate_185(n336,n330,n335);
and gate_186(n337,pi26,n185);
not gate_187(n338,n337);
and gate_188(n339,pi30,n186);
not gate_189(n340,n339);
and gate_190(n341,n338,n340);
not gate_191(n342,n341);
and gate_192(n343,n228,n342);
not gate_193(n344,n343);
and gate_194(n345,n336,n344);
not gate_195(po06,n345);
and gate_196(n347,pi24,n218);
not gate_197(n348,n347);
and gate_198(n349,pi16,n185);
not gate_199(n350,n349);
and gate_200(n351,n217,n349);
not gate_201(n352,n351);
and gate_202(n353,n214,n352);
and gate_203(n354,n348,n353);
and gate_204(n355,pi27,n185);
not gate_205(n356,n355);
and gate_206(n357,pi31,n186);
not gate_207(n358,n357);
and gate_208(n359,n356,n358);
not gate_209(n360,n359);
and gate_210(n361,n228,n360);
not gate_211(n362,n361);
and gate_212(n363,n354,n362);
not gate_213(po07,n363);
and gate_214(n365,pi25,n218);
not gate_215(n366,n365);
and gate_216(n367,pi17,n185);
not gate_217(n368,n367);
and gate_218(n369,n217,n367);
not gate_219(n370,n369);
and gate_220(n371,n214,n370);
and gate_221(n372,n366,n371);
and gate_222(n373,pi28,n185);
not gate_223(n374,n373);
and gate_224(n375,pi32,n186);
not gate_225(n376,n375);
and gate_226(n377,n374,n376);
not gate_227(n378,n377);
and gate_228(n379,n228,n378);
not gate_229(n380,n379);
and gate_230(n381,n372,n380);
not gate_231(po08,n381);
and gate_232(n383,pi26,n218);
not gate_233(n384,n383);
and gate_234(n385,pi18,n185);
not gate_235(n386,n385);
and gate_236(n387,n217,n385);
not gate_237(n388,n387);
and gate_238(n389,n214,n388);
and gate_239(n390,n384,n389);
and gate_240(n391,pi29,n185);
not gate_241(n392,n391);
and gate_242(n393,pi33,n186);
not gate_243(n394,n393);
and gate_244(n395,n392,n394);
not gate_245(n396,n395);
and gate_246(n397,n228,n396);
not gate_247(n398,n397);
and gate_248(n399,n390,n398);
not gate_249(po09,n399);
and gate_250(n401,pi27,n218);
not gate_251(n402,n401);
and gate_252(n403,pi19,n185);
not gate_253(n404,n403);
and gate_254(n405,n217,n403);
not gate_255(n406,n405);
and gate_256(n407,n214,n406);
and gate_257(n408,n402,n407);
and gate_258(n409,pi30,n185);
not gate_259(n410,n409);
and gate_260(n411,pi34,n186);
not gate_261(n412,n411);
and gate_262(n413,n410,n412);
not gate_263(n414,n413);
and gate_264(n415,n228,n414);
not gate_265(n416,n415);
and gate_266(n417,n408,n416);
not gate_267(po10,n417);
and gate_268(n419,pi28,n218);
not gate_269(n420,n419);
and gate_270(n421,n217,n229);
not gate_271(n422,n421);
and gate_272(n423,n214,n422);
and gate_273(n424,n420,n423);
and gate_274(n425,pi31,n185);
not gate_275(n426,n425);
and gate_276(n427,pi35,n186);
not gate_277(n428,n427);
and gate_278(n429,n426,n428);
not gate_279(n430,n429);
and gate_280(n431,n228,n430);
not gate_281(n432,n431);
and gate_282(n433,n424,n432);
not gate_283(po11,n433);
and gate_284(n435,pi29,n218);
not gate_285(n436,n435);
and gate_286(n437,n217,n247);
not gate_287(n438,n437);
and gate_288(n439,n214,n438);
and gate_289(n440,n436,n439);
and gate_290(n441,pi32,n185);
not gate_291(n442,n441);
and gate_292(n443,pi36,n186);
not gate_293(n444,n443);
and gate_294(n445,n442,n444);
not gate_295(n446,n445);
and gate_296(n447,n228,n446);
not gate_297(n448,n447);
and gate_298(n449,n440,n448);
not gate_299(po12,n449);
and gate_300(n451,pi30,n218);
not gate_301(n452,n451);
and gate_302(n453,n217,n265);
not gate_303(n454,n453);
and gate_304(n455,n214,n454);
and gate_305(n456,n452,n455);
and gate_306(n457,pi33,n185);
not gate_307(n458,n457);
and gate_308(n459,pi37,n186);
not gate_309(n460,n459);
and gate_310(n461,n458,n460);
not gate_311(n462,n461);
and gate_312(n463,n228,n462);
not gate_313(n464,n463);
and gate_314(n465,n456,n464);
not gate_315(po13,n465);
and gate_316(n467,pi31,n218);
not gate_317(n468,n467);
and gate_318(n469,n217,n283);
not gate_319(n470,n469);
and gate_320(n471,n214,n470);
and gate_321(n472,n468,n471);
and gate_322(n473,pi34,n185);
not gate_323(n474,n473);
and gate_324(n475,pi38,n186);
not gate_325(n476,n475);
and gate_326(n477,n474,n476);
not gate_327(n478,n477);
and gate_328(n479,n228,n478);
not gate_329(n480,n479);
and gate_330(n481,n472,n480);
not gate_331(po14,n481);
and gate_332(n483,pi32,n218);
not gate_333(n484,n483);
and gate_334(n485,n217,n301);
not gate_335(n486,n485);
and gate_336(n487,n214,n486);
and gate_337(n488,n484,n487);
and gate_338(n489,pi35,n185);
not gate_339(n490,n489);
and gate_340(n491,pi39,n186);
not gate_341(n492,n491);
and gate_342(n493,n490,n492);
not gate_343(n494,n493);
and gate_344(n495,n228,n494);
not gate_345(n496,n495);
and gate_346(n497,n488,n496);
not gate_347(po15,n497);
and gate_348(n499,pi33,n218);
not gate_349(n500,n499);
and gate_350(n501,n217,n319);
not gate_351(n502,n501);
and gate_352(n503,n214,n502);
and gate_353(n504,n500,n503);
and gate_354(n505,pi36,n185);
not gate_355(n506,n505);
and gate_356(n507,pi52,n186);
not gate_357(n508,n507);
and gate_358(n509,n506,n508);
not gate_359(n510,n509);
and gate_360(n511,n228,n510);
not gate_361(n512,n511);
and gate_362(n513,n504,n512);
not gate_363(po16,n513);
and gate_364(n515,pi34,n218);
not gate_365(n516,n515);
and gate_366(n517,n217,n337);
not gate_367(n518,n517);
and gate_368(n519,n214,n518);
and gate_369(n520,n516,n519);
and gate_370(n521,pi37,n185);
not gate_371(n522,n521);
and gate_372(n523,pi53,n186);
not gate_373(n524,n523);
and gate_374(n525,n522,n524);
not gate_375(n526,n525);
and gate_376(n527,n228,n526);
not gate_377(n528,n527);
and gate_378(n529,n520,n528);
not gate_379(po17,n529);
and gate_380(n531,pi35,n218);
not gate_381(n532,n531);
and gate_382(n533,n217,n355);
not gate_383(n534,n533);
and gate_384(n535,n214,n534);
and gate_385(n536,n532,n535);
and gate_386(n537,pi38,n185);
not gate_387(n538,n537);
and gate_388(n539,pi54,n186);
not gate_389(n540,n539);
and gate_390(n541,n538,n540);
not gate_391(n542,n541);
and gate_392(n543,n228,n542);
not gate_393(n544,n543);
and gate_394(n545,n536,n544);
not gate_395(po18,n545);
and gate_396(n547,pi36,n218);
not gate_397(n548,n547);
and gate_398(n549,n217,n373);
not gate_399(n550,n549);
and gate_400(n551,n214,n550);
and gate_401(n552,n548,n551);
and gate_402(n553,pi39,n185);
not gate_403(n554,n553);
and gate_404(n555,pi55,n186);
not gate_405(n556,n555);
and gate_406(n557,n554,n556);
not gate_407(n558,n557);
and gate_408(n559,n228,n558);
not gate_409(n560,n559);
and gate_410(n561,n552,n560);
not gate_411(po19,n561);
and gate_412(n563,pi41,n185);
not gate_413(n564,n563);
and gate_414(n565,n228,n563);
not gate_415(n566,n565);
and gate_416(n567,pi56,n186);
and gate_417(n568,n228,n567);
not gate_418(n569,n568);
and gate_419(n570,n566,n569);
and gate_420(n571,pi37,n218);
not gate_421(n572,n571);
and gate_422(n573,n217,n391);
not gate_423(n574,n573);
and gate_424(n575,n214,n574);
and gate_425(n576,n572,n575);
and gate_426(n577,n570,n576);
not gate_427(po20,n577);
and gate_428(n579,pi42,n185);
not gate_429(n580,n579);
and gate_430(n581,n228,n579);
not gate_431(n582,n581);
and gate_432(n583,pi57,n186);
and gate_433(n584,n228,n583);
not gate_434(n585,n584);
and gate_435(n586,n582,n585);
and gate_436(n587,pi38,n218);
not gate_437(n588,n587);
and gate_438(n589,n217,n409);
not gate_439(n590,n589);
and gate_440(n591,n214,n590);
and gate_441(n592,n588,n591);
and gate_442(n593,n586,n592);
not gate_443(po21,n593);
and gate_444(n595,pi43,n185);
not gate_445(n596,n595);
and gate_446(n597,n228,n595);
not gate_447(n598,n597);
and gate_448(n599,pi58,n186);
and gate_449(n600,n228,n599);
not gate_450(n601,n600);
and gate_451(n602,n598,n601);
and gate_452(n603,pi39,n218);
not gate_453(n604,n603);
and gate_454(n605,n217,n425);
not gate_455(n606,n605);
and gate_456(n607,n214,n606);
and gate_457(n608,n604,n607);
and gate_458(n609,n602,n608);
not gate_459(po22,n609);
and gate_460(n611,pi44,n185);
not gate_461(n612,n611);
and gate_462(n613,n228,n611);
not gate_463(n614,n613);
and gate_464(n615,pi59,n186);
and gate_465(n616,n228,n615);
not gate_466(n617,n616);
and gate_467(n618,n614,n617);
and gate_468(n619,pi40,n218);
not gate_469(n620,n619);
and gate_470(n621,n217,n441);
not gate_471(n622,n621);
and gate_472(n623,n214,n622);
and gate_473(n624,n620,n623);
and gate_474(n625,n618,n624);
not gate_475(po23,n625);
and gate_476(n627,pi45,n185);
not gate_477(n628,n627);
and gate_478(n629,n228,n627);
not gate_479(n630,n629);
and gate_480(n631,pi60,n186);
and gate_481(n632,n228,n631);
not gate_482(n633,n632);
and gate_483(n634,n630,n633);
and gate_484(n635,n217,n457);
not gate_485(n636,n635);
and gate_486(n637,n214,n636);
and gate_487(n638,n219,n637);
and gate_488(n639,n634,n638);
not gate_489(po24,n639);
and gate_490(n641,pi46,n185);
not gate_491(n642,n641);
and gate_492(n643,n228,n641);
not gate_493(n644,n643);
and gate_494(n645,pi61,n186);
and gate_495(n646,n228,n645);
not gate_496(n647,n646);
and gate_497(n648,n644,n647);
and gate_498(n649,n217,n473);
not gate_499(n650,n649);
and gate_500(n651,n214,n650);
and gate_501(n652,n219,n651);
and gate_502(n653,n648,n652);
not gate_503(po25,n653);
and gate_504(n655,pi47,n185);
not gate_505(n656,n655);
and gate_506(n657,n228,n655);
not gate_507(n658,n657);
and gate_508(n659,pi62,n186);
and gate_509(n660,n228,n659);
not gate_510(n661,n660);
and gate_511(n662,n658,n661);
and gate_512(n663,n217,n489);
not gate_513(n664,n663);
and gate_514(n665,n214,n664);
and gate_515(n666,n219,n665);
and gate_516(n667,n662,n666);
not gate_517(po26,n667);
and gate_518(n669,pi48,n185);
not gate_519(n670,n669);
and gate_520(n671,n228,n669);
not gate_521(n672,n671);
and gate_522(n673,pi63,n186);
and gate_523(n674,n228,n673);
not gate_524(n675,n674);
and gate_525(n676,n672,n675);
and gate_526(n677,n217,n505);
not gate_527(n678,n677);
and gate_528(n679,n214,n678);
and gate_529(n680,n219,n679);
and gate_530(n681,n676,n680);
not gate_531(po27,n681);
and gate_532(n683,pi49,n185);
not gate_533(n684,n683);
and gate_534(n685,n228,n683);
not gate_535(n686,n685);
and gate_536(n687,pi64,n186);
and gate_537(n688,n228,n687);
not gate_538(n689,n688);
and gate_539(n690,n686,n689);
and gate_540(n691,n217,n521);
not gate_541(n692,n691);
and gate_542(n693,n214,n692);
and gate_543(n694,n219,n693);
and gate_544(n695,n690,n694);
not gate_545(po28,n695);
and gate_546(n697,pi50,n185);
not gate_547(n698,n697);
and gate_548(n699,n228,n697);
not gate_549(n700,n699);
and gate_550(n701,pi65,n186);
and gate_551(n702,n228,n701);
not gate_552(n703,n702);
and gate_553(n704,n700,n703);
and gate_554(n705,n217,n537);
not gate_555(n706,n705);
and gate_556(n707,n214,n706);
and gate_557(n708,n219,n707);
and gate_558(n709,n704,n708);
not gate_559(po29,n709);
and gate_560(n711,pi51,n185);
not gate_561(n712,n711);
and gate_562(n713,n228,n711);
not gate_563(n714,n713);
and gate_564(n715,pi66,n186);
and gate_565(n716,n228,n715);
not gate_566(n717,n716);
and gate_567(n718,n714,n717);
and gate_568(n719,n217,n553);
not gate_569(n720,n719);
and gate_570(n721,n214,n720);
and gate_571(n722,n219,n721);
and gate_572(n723,n718,n722);
not gate_573(po30,n723);
and gate_574(n725,pi87,n186);
not gate_575(n726,n725);
and gate_576(n727,n228,n725);
not gate_577(n728,n727);
and gate_578(n729,n672,n728);
and gate_579(n730,pi83,n185);
not gate_580(n731,n730);
and gate_581(n732,pi45,n186);
not gate_582(n733,n732);
and gate_583(n734,n731,n733);
not gate_584(n735,n734);
and gate_585(n736,n217,n735);
not gate_586(n737,n736);
and gate_587(n738,n729,n737);
and gate_588(n739,n214,n738);
not gate_589(po31,n739);
and gate_590(n741,pi09,n186);
not gate_591(n742,n741);
and gate_592(n743,n228,n741);
not gate_593(n744,n743);
and gate_594(n745,n686,n744);
and gate_595(n746,pi84,n185);
not gate_596(n747,n746);
and gate_597(n748,pi46,n186);
not gate_598(n749,n748);
and gate_599(n750,n747,n749);
not gate_600(n751,n750);
and gate_601(n752,n217,n751);
not gate_602(n753,n752);
and gate_603(n754,n745,n753);
and gate_604(n755,n214,n754);
not gate_605(po32,n755);
and gate_606(n757,pi10,n186);
not gate_607(n758,n757);
and gate_608(n759,n228,n757);
not gate_609(n760,n759);
and gate_610(n761,n700,n760);
and gate_611(n762,pi85,n185);
not gate_612(n763,n762);
and gate_613(n764,pi47,n186);
not gate_614(n765,n764);
and gate_615(n766,n763,n765);
not gate_616(n767,n766);
and gate_617(n768,n217,n767);
not gate_618(n769,n768);
and gate_619(n770,n761,n769);
and gate_620(n771,n214,n770);
not gate_621(po33,n771);
and gate_622(n773,pi11,n186);
not gate_623(n774,n773);
and gate_624(n775,n228,n773);
not gate_625(n776,n775);
and gate_626(n777,n714,n776);
and gate_627(n778,pi86,n185);
not gate_628(n779,n778);
and gate_629(n780,pi48,n186);
not gate_630(n781,n780);
and gate_631(n782,n779,n781);
not gate_632(n783,n782);
and gate_633(n784,n217,n783);
not gate_634(n785,n784);
and gate_635(n786,n777,n785);
and gate_636(n787,n214,n786);
not gate_637(po34,n787);
and gate_638(n789,pi49,n186);
not gate_639(n790,n789);
and gate_640(n791,n564,n790);
not gate_641(n792,n791);
and gate_642(n793,n217,n792);
not gate_643(n794,n793);
and gate_644(n795,pi87,n185);
not gate_645(n796,n795);
and gate_646(n797,pi12,n186);
not gate_647(n798,n797);
and gate_648(n799,n796,n798);
not gate_649(n800,n799);
and gate_650(n801,n228,n800);
not gate_651(n802,n801);
and gate_652(n803,n794,n802);
and gate_653(n804,n214,n803);
not gate_654(po35,n804);
and gate_655(n806,pi50,n186);
not gate_656(n807,n806);
and gate_657(n808,n580,n807);
not gate_658(n809,n808);
and gate_659(n810,n217,n809);
not gate_660(n811,n810);
and gate_661(n812,pi13,n186);
not gate_662(n813,n812);
and gate_663(n814,n223,n813);
not gate_664(n815,n814);
and gate_665(n816,n228,n815);
not gate_666(n817,n816);
and gate_667(n818,n811,n817);
and gate_668(n819,n214,n818);
not gate_669(po36,n819);
and gate_670(n821,pi51,n186);
not gate_671(n822,n821);
and gate_672(n823,n596,n822);
not gate_673(n824,n823);
and gate_674(n825,n217,n824);
not gate_675(n826,n825);
and gate_676(n827,pi14,n186);
not gate_677(n828,n827);
and gate_678(n829,n242,n828);
not gate_679(n830,n829);
and gate_680(n831,n228,n830);
not gate_681(n832,n831);
and gate_682(n833,n826,n832);
and gate_683(n834,n214,n833);
not gate_684(po37,n834);
and gate_685(n836,n612,n726);
not gate_686(n837,n836);
and gate_687(n838,n217,n837);
not gate_688(n839,n838);
and gate_689(n840,pi15,n186);
not gate_690(n841,n840);
and gate_691(n842,n260,n841);
not gate_692(n843,n842);
and gate_693(n844,n228,n843);
not gate_694(n845,n844);
and gate_695(n846,n839,n845);
and gate_696(n847,n214,n846);
not gate_697(po38,n847);
and gate_698(n849,n628,n742);
not gate_699(n850,n849);
and gate_700(n851,n217,n850);
not gate_701(n852,n851);
and gate_702(n853,pi16,n186);
not gate_703(n854,n853);
and gate_704(n855,n278,n854);
not gate_705(n856,n855);
and gate_706(n857,n228,n856);
not gate_707(n858,n857);
and gate_708(n859,n852,n858);
and gate_709(n860,n214,n859);
not gate_710(po39,n860);
and gate_711(n862,n642,n758);
not gate_712(n863,n862);
and gate_713(n864,n217,n863);
not gate_714(n865,n864);
and gate_715(n866,pi17,n186);
not gate_716(n867,n866);
and gate_717(n868,n296,n867);
not gate_718(n869,n868);
and gate_719(n870,n228,n869);
not gate_720(n871,n870);
and gate_721(n872,n865,n871);
and gate_722(n873,n214,n872);
not gate_723(po40,n873);
and gate_724(n875,n656,n774);
not gate_725(n876,n875);
and gate_726(n877,n217,n876);
not gate_727(n878,n877);
and gate_728(n879,pi18,n186);
not gate_729(n880,n879);
and gate_730(n881,n314,n880);
not gate_731(n882,n881);
and gate_732(n883,n228,n882);
not gate_733(n884,n883);
and gate_734(n885,n878,n884);
and gate_735(n886,n214,n885);
not gate_736(po41,n886);
and gate_737(n888,n670,n798);
not gate_738(n889,n888);
and gate_739(n890,n217,n889);
not gate_740(n891,n890);
and gate_741(n892,pi19,n186);
not gate_742(n893,n892);
and gate_743(n894,n332,n893);
not gate_744(n895,n894);
and gate_745(n896,n228,n895);
not gate_746(n897,n896);
and gate_747(n898,n891,n897);
and gate_748(n899,n214,n898);
not gate_749(po42,n899);
and gate_750(n901,n684,n813);
not gate_751(n902,n901);
and gate_752(n903,n217,n902);
not gate_753(n904,n903);
and gate_754(n905,pi20,n186);
not gate_755(n906,n905);
and gate_756(n907,n350,n906);
not gate_757(n908,n907);
and gate_758(n909,n228,n908);
not gate_759(n910,n909);
and gate_760(n911,n904,n910);
and gate_761(n912,n214,n911);
not gate_762(po43,n912);
and gate_763(n914,n698,n828);
not gate_764(n915,n914);
and gate_765(n916,n217,n915);
not gate_766(n917,n916);
and gate_767(n918,pi21,n186);
not gate_768(n919,n918);
and gate_769(n920,n368,n919);
not gate_770(n921,n920);
and gate_771(n922,n228,n921);
not gate_772(n923,n922);
and gate_773(n924,n917,n923);
and gate_774(n925,n214,n924);
not gate_775(po44,n925);
and gate_776(n927,n712,n841);
not gate_777(n928,n927);
and gate_778(n929,n217,n928);
not gate_779(n930,n929);
and gate_780(n931,pi22,n186);
not gate_781(n932,n931);
and gate_782(n933,n386,n932);
not gate_783(n934,n933);
and gate_784(n935,n228,n934);
not gate_785(n936,n935);
and gate_786(n937,n930,n936);
and gate_787(n938,n214,n937);
not gate_788(po45,n938);
and gate_789(n940,n796,n854);
not gate_790(n941,n940);
and gate_791(n942,n217,n941);
not gate_792(n943,n942);
and gate_793(n944,pi23,n186);
not gate_794(n945,n944);
and gate_795(n946,n404,n945);
not gate_796(n947,n946);
and gate_797(n948,n228,n947);
not gate_798(n949,n948);
and gate_799(n950,n943,n949);
and gate_800(n951,n214,n950);
not gate_801(po46,n951);
and gate_802(n953,pi67,n185);
not gate_803(n954,n953);
and gate_804(n955,pi75,n186);
not gate_805(n956,n955);
and gate_806(n957,n954,n956);
not gate_807(n958,n957);
and gate_808(n959,n217,n958);
not gate_809(n960,n959);
and gate_810(n961,pi78,n185);
not gate_811(n962,n961);
and gate_812(n963,pi82,n186);
not gate_813(n964,n963);
and gate_814(n965,n962,n964);
not gate_815(n966,n965);
and gate_816(n967,n228,n966);
not gate_817(n968,n967);
and gate_818(n969,n960,n968);
and gate_819(n970,n214,n969);
not gate_820(po47,n970);
and gate_821(n972,pi68,n185);
not gate_822(n973,n972);
and gate_823(n974,pi76,n186);
not gate_824(n975,n974);
and gate_825(n976,n973,n975);
not gate_826(n977,n976);
and gate_827(n978,n217,n977);
not gate_828(n979,n978);
and gate_829(n980,pi79,n185);
not gate_830(n981,n980);
and gate_831(n982,pi83,n186);
not gate_832(n983,n982);
and gate_833(n984,n981,n983);
not gate_834(n985,n984);
and gate_835(n986,n228,n985);
not gate_836(n987,n986);
and gate_837(n988,n979,n987);
and gate_838(n989,n214,n988);
not gate_839(po48,n989);
and gate_840(n991,pi69,n185);
not gate_841(n992,n991);
and gate_842(n993,pi77,n186);
not gate_843(n994,n993);
and gate_844(n995,n992,n994);
not gate_845(n996,n995);
and gate_846(n997,n217,n996);
not gate_847(n998,n997);
and gate_848(n999,pi80,n185);
not gate_849(n1000,n999);
and gate_850(n1001,pi84,n186);
not gate_851(n1002,n1001);
and gate_852(n1003,n1000,n1002);
not gate_853(n1004,n1003);
and gate_854(n1005,n228,n1004);
not gate_855(n1006,n1005);
and gate_856(n1007,n998,n1006);
and gate_857(n1008,n214,n1007);
not gate_858(po49,n1008);
and gate_859(n1010,pi70,n185);
not gate_860(n1011,n1010);
and gate_861(n1012,pi78,n186);
not gate_862(n1013,n1012);
and gate_863(n1014,n1011,n1013);
not gate_864(n1015,n1014);
and gate_865(n1016,n217,n1015);
not gate_866(n1017,n1016);
and gate_867(n1018,pi81,n185);
not gate_868(n1019,n1018);
and gate_869(n1020,pi85,n186);
not gate_870(n1021,n1020);
and gate_871(n1022,n1019,n1021);
not gate_872(n1023,n1022);
and gate_873(n1024,n228,n1023);
not gate_874(n1025,n1024);
and gate_875(n1026,n1017,n1025);
and gate_876(n1027,n214,n1026);
not gate_877(po50,n1027);
and gate_878(n1029,pi71,n185);
not gate_879(n1030,n1029);
and gate_880(n1031,pi79,n186);
not gate_881(n1032,n1031);
and gate_882(n1033,n1030,n1032);
not gate_883(n1034,n1033);
and gate_884(n1035,n217,n1034);
not gate_885(n1036,n1035);
and gate_886(n1037,pi82,n185);
not gate_887(n1038,n1037);
and gate_888(n1039,pi86,n186);
not gate_889(n1040,n1039);
and gate_890(n1041,n1038,n1040);
not gate_891(n1042,n1041);
and gate_892(n1043,n228,n1042);
not gate_893(n1044,n1043);
and gate_894(n1045,n1036,n1044);
and gate_895(n1046,n214,n1045);
not gate_896(po51,n1046);
and gate_897(n1048,pi72,n185);
not gate_898(n1049,n1048);
and gate_899(n1050,pi80,n186);
not gate_900(n1051,n1050);
and gate_901(n1052,n1049,n1051);
not gate_902(n1053,n1052);
and gate_903(n1054,n217,n1053);
not gate_904(n1055,n1054);
and gate_905(n1056,pi41,n186);
not gate_906(n1057,n1056);
and gate_907(n1058,n731,n1057);
not gate_908(n1059,n1058);
and gate_909(n1060,n228,n1059);
not gate_910(n1061,n1060);
and gate_911(n1062,n1055,n1061);
and gate_912(n1063,n214,n1062);
not gate_913(po52,n1063);
and gate_914(n1065,pi73,n185);
not gate_915(n1066,n1065);
and gate_916(n1067,pi81,n186);
not gate_917(n1068,n1067);
and gate_918(n1069,n1066,n1068);
not gate_919(n1070,n1069);
and gate_920(n1071,n217,n1070);
not gate_921(n1072,n1071);
and gate_922(n1073,pi42,n186);
not gate_923(n1074,n1073);
and gate_924(n1075,n747,n1074);
not gate_925(n1076,n1075);
and gate_926(n1077,n228,n1076);
not gate_927(n1078,n1077);
and gate_928(n1079,n1072,n1078);
and gate_929(n1080,n214,n1079);
not gate_930(po53,n1080);
and gate_931(n1082,pi74,n185);
not gate_932(n1083,n1082);
and gate_933(n1084,n964,n1083);
not gate_934(n1085,n1084);
and gate_935(n1086,n217,n1085);
not gate_936(n1087,n1086);
and gate_937(n1088,pi43,n186);
not gate_938(n1089,n1088);
and gate_939(n1090,n763,n1089);
not gate_940(n1091,n1090);
and gate_941(n1092,n228,n1091);
not gate_942(n1093,n1092);
and gate_943(n1094,n1087,n1093);
and gate_944(n1095,n214,n1094);
not gate_945(po54,n1095);
and gate_946(n1097,pi75,n185);
not gate_947(n1098,n1097);
and gate_948(n1099,n983,n1098);
not gate_949(n1100,n1099);
and gate_950(n1101,n217,n1100);
not gate_951(n1102,n1101);
and gate_952(n1103,pi44,n186);
not gate_953(n1104,n1103);
and gate_954(n1105,n779,n1104);
not gate_955(n1106,n1105);
and gate_956(n1107,n228,n1106);
not gate_957(n1108,n1107);
and gate_958(n1109,n1102,n1108);
and gate_959(n1110,n214,n1109);
not gate_960(po55,n1110);
and gate_961(n1112,n228,n732);
not gate_962(n1113,n1112);
and gate_963(n1114,n566,n1113);
and gate_964(n1115,pi76,n185);
not gate_965(n1116,n1115);
and gate_966(n1117,n1002,n1116);
not gate_967(n1118,n1117);
and gate_968(n1119,n217,n1118);
not gate_969(n1120,n1119);
and gate_970(n1121,n1114,n1120);
and gate_971(n1122,n214,n1121);
not gate_972(po56,n1122);
and gate_973(n1124,n228,n748);
not gate_974(n1125,n1124);
and gate_975(n1126,n582,n1125);
and gate_976(n1127,pi77,n185);
not gate_977(n1128,n1127);
and gate_978(n1129,n1021,n1128);
not gate_979(n1130,n1129);
and gate_980(n1131,n217,n1130);
not gate_981(n1132,n1131);
and gate_982(n1133,n1126,n1132);
and gate_983(n1134,n214,n1133);
not gate_984(po57,n1134);
and gate_985(n1136,n228,n764);
not gate_986(n1137,n1136);
and gate_987(n1138,n598,n1137);
and gate_988(n1139,n962,n1040);
not gate_989(n1140,n1139);
and gate_990(n1141,n217,n1140);
not gate_991(n1142,n1141);
and gate_992(n1143,n1138,n1142);
and gate_993(n1144,n214,n1143);
not gate_994(po58,n1144);
and gate_995(n1146,n228,n780);
not gate_996(n1147,n1146);
and gate_997(n1148,n614,n1147);
and gate_998(n1149,n981,n1057);
not gate_999(n1150,n1149);
and gate_1000(n1151,n217,n1150);
not gate_1001(n1152,n1151);
and gate_1002(n1153,n1148,n1152);
and gate_1003(n1154,n214,n1153);
not gate_1004(po59,n1154);
and gate_1005(n1156,n228,n789);
not gate_1006(n1157,n1156);
and gate_1007(n1158,n630,n1157);
and gate_1008(n1159,n1000,n1074);
not gate_1009(n1160,n1159);
and gate_1010(n1161,n217,n1160);
not gate_1011(n1162,n1161);
and gate_1012(n1163,n1158,n1162);
and gate_1013(n1164,n214,n1163);
not gate_1014(po60,n1164);
and gate_1015(n1166,n228,n806);
not gate_1016(n1167,n1166);
and gate_1017(n1168,n644,n1167);
and gate_1018(n1169,n1019,n1089);
not gate_1019(n1170,n1169);
and gate_1020(n1171,n217,n1170);
not gate_1021(n1172,n1171);
and gate_1022(n1173,n1168,n1172);
and gate_1023(n1174,n214,n1173);
not gate_1024(po61,n1174);
and gate_1025(n1176,n228,n821);
not gate_1026(n1177,n1176);
and gate_1027(n1178,n658,n1177);
and gate_1028(n1179,n1038,n1104);
not gate_1029(n1180,n1179);
and gate_1030(n1181,n217,n1180);
not gate_1031(n1182,n1181);
and gate_1032(n1183,n1178,n1182);
and gate_1033(n1184,n214,n1183);
not gate_1034(po62,n1184);
endmodule
