// Verilog File 
module c432 (G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat,G223gat,G329gat,G370gat,
G421gat,G430gat,G431gat,G432gat);

input G1gat,G4gat,G8gat,G11gat,G14gat,G17gat,G21gat,G24gat,G27gat,
G30gat,G34gat,G37gat,G40gat,G43gat,G47gat,G50gat,G53gat,G56gat,G60gat,
G63gat,G66gat,G69gat,G73gat,G76gat,G79gat,G82gat,G86gat,G89gat,G92gat,
G95gat,G99gat,G102gat,G105gat,G108gat,G112gat,G115gat;

output G223gat,G329gat,G370gat,G421gat,G430gat,G431gat,G432gat;

wire G118gat,G119gat,G122gat,G123gat,G126gat,G127gat,G130gat,G131gat,G134gat,
G135gat,G138gat,G139gat,G142gat,G143gat,G146gat,G147gat,G150gat,G151gat,G154gat,
G157gat,G158gat,G159gat,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat,
G183gat,G184gat,G185gat,G186gat,G187gat,G188gat,G189gat,G190gat,G191gat,G192gat,
G193gat,G194gat,G195gat,G196gat,G197gat,G198gat,G199gat,G203gat,G213gat,G224gat,
G227gat,G230gat,G233gat,G236gat,G239gat,G242gat,G243gat,G246gat,G247gat,G250gat,
G251gat,G254gat,G255gat,G256gat,G257gat,G258gat,G259gat,G260gat,G263gat,G264gat,
G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat,G288gat,G289gat,G290gat,
G291gat,G292gat,G293gat,G294gat,G295gat,G296gat,G300gat,G301gat,G302gat,G303gat,
G304gat,G305gat,G306gat,G307gat,G308gat,G309gat,G319gat,G330gat,G331gat,G332gat,
G333gat,G334gat,G335gat,G336gat,G337gat,G338gat,G339gat,G340gat,G341gat,G342gat,
G343gat,G344gat,G345gat,G346gat,G347gat,G348gat,G349gat,G350gat,G351gat,G352gat,
G353gat,G354gat,G355gat,G356gat,G357gat,G360gat,G371gat,G372gat,G373gat,G374gat,
G375gat,G376gat,G377gat,G378gat,G379gat,G380gat,G381gat,G386gat,G393gat,G399gat,
G404gat,G407gat,G411gat,G414gat,G415gat,G416gat,G417gat,G418gat,G419gat,G420gat,
G422gat,G425gat,G428gat,G429gat;
not gate_0(G118gat,G1gat);
not gate_1(G119gat,G4gat);
not gate_2(G122gat,G11gat);
not gate_3(G123gat,G17gat);
not gate_4(G126gat,G24gat);
not gate_5(G127gat,G30gat);
not gate_6(G130gat,G37gat);
not gate_7(G131gat,G43gat);
not gate_8(G134gat,G50gat);
not gate_9(G135gat,G56gat);
not gate_10(G138gat,G63gat);
not gate_11(G139gat,G69gat);
not gate_12(G142gat,G76gat);
not gate_13(G143gat,G82gat);
not gate_14(G146gat,G89gat);
not gate_15(G147gat,G95gat);
not gate_16(G150gat,G102gat);
not gate_17(G151gat,G108gat);
nand gate_18(G154gat,G118gat,G4gat);
nor gate_19(G157gat,G8gat,G119gat);
nor gate_20(G158gat,G14gat,G119gat);
nand gate_21(G159gat,G122gat,G17gat);
nand gate_22(G162gat,G126gat,G30gat);
nand gate_23(G165gat,G130gat,G43gat);
nand gate_24(G168gat,G134gat,G56gat);
nand gate_25(G171gat,G138gat,G69gat);
nand gate_26(G174gat,G142gat,G82gat);
nand gate_27(G177gat,G146gat,G95gat);
nand gate_28(G180gat,G150gat,G108gat);
nor gate_29(G183gat,G21gat,G123gat);
nor gate_30(G184gat,G27gat,G123gat);
nor gate_31(G185gat,G34gat,G127gat);
nor gate_32(G186gat,G40gat,G127gat);
nor gate_33(G187gat,G47gat,G131gat);
nor gate_34(G188gat,G53gat,G131gat);
nor gate_35(G189gat,G60gat,G135gat);
nor gate_36(G190gat,G66gat,G135gat);
nor gate_37(G191gat,G73gat,G139gat);
nor gate_38(G192gat,G79gat,G139gat);
nor gate_39(G193gat,G86gat,G143gat);
nor gate_40(G194gat,G92gat,G143gat);
nor gate_41(G195gat,G99gat,G147gat);
nor gate_42(G196gat,G105gat,G147gat);
nor gate_43(G197gat,G112gat,G151gat);
nor gate_44(G198gat,G115gat,G151gat);
and gate_45(G199gat,G154gat,G159gat,G162gat,G165gat,G168gat,G171gat,G174gat,G177gat,G180gat);
not gate_46(G203gat,G199gat);
not gate_47(G213gat,G199gat);
not gate_48(G223gat,G199gat);
xor gate_49(G224gat,G203gat,G154gat);
xor gate_50(G227gat,G203gat,G159gat);
xor gate_51(G230gat,G203gat,G162gat);
xor gate_52(G233gat,G203gat,G165gat);
xor gate_53(G236gat,G203gat,G168gat);
xor gate_54(G239gat,G203gat,G171gat);
nand gate_55(G242gat,G1gat,G213gat);
xor gate_56(G243gat,G203gat,G174gat);
nand gate_57(G246gat,G213gat,G11gat);
xor gate_58(G247gat,G203gat,G177gat);
nand gate_59(G250gat,G213gat,G24gat);
xor gate_60(G251gat,G203gat,G180gat);
nand gate_61(G254gat,G213gat,G37gat);
nand gate_62(G255gat,G213gat,G50gat);
nand gate_63(G256gat,G213gat,G63gat);
nand gate_64(G257gat,G213gat,G76gat);
nand gate_65(G258gat,G213gat,G89gat);
nand gate_66(G259gat,G213gat,G102gat);
nand gate_67(G260gat,G224gat,G157gat);
nand gate_68(G263gat,G224gat,G158gat);
nand gate_69(G264gat,G227gat,G183gat);
nand gate_70(G267gat,G230gat,G185gat);
nand gate_71(G270gat,G233gat,G187gat);
nand gate_72(G273gat,G236gat,G189gat);
nand gate_73(G276gat,G239gat,G191gat);
nand gate_74(G279gat,G243gat,G193gat);
nand gate_75(G282gat,G247gat,G195gat);
nand gate_76(G285gat,G251gat,G197gat);
nand gate_77(G288gat,G227gat,G184gat);
nand gate_78(G289gat,G230gat,G186gat);
nand gate_79(G290gat,G233gat,G188gat);
nand gate_80(G291gat,G236gat,G190gat);
nand gate_81(G292gat,G239gat,G192gat);
nand gate_82(G293gat,G243gat,G194gat);
nand gate_83(G294gat,G247gat,G196gat);
nand gate_84(G295gat,G251gat,G198gat);
and gate_85(G296gat,G260gat,G264gat,G267gat,G270gat,G273gat,G276gat,G279gat,G282gat,G285gat);
not gate_86(G300gat,G263gat);
not gate_87(G301gat,G288gat);
not gate_88(G302gat,G289gat);
not gate_89(G303gat,G290gat);
not gate_90(G304gat,G291gat);
not gate_91(G305gat,G292gat);
not gate_92(G306gat,G293gat);
not gate_93(G307gat,G294gat);
not gate_94(G308gat,G295gat);
not gate_95(G309gat,G296gat);
not gate_96(G319gat,G296gat);
not gate_97(G329gat,G296gat);
xor gate_98(G330gat,G309gat,G260gat);
xor gate_99(G331gat,G309gat,G264gat);
xor gate_100(G332gat,G309gat,G267gat);
xor gate_101(G333gat,G309gat,G270gat);
nand gate_102(G334gat,G8gat,G319gat);
xor gate_103(G335gat,G309gat,G273gat);
nand gate_104(G336gat,G319gat,G21gat);
xor gate_105(G337gat,G309gat,G276gat);
nand gate_106(G338gat,G319gat,G34gat);
xor gate_107(G339gat,G309gat,G279gat);
nand gate_108(G340gat,G319gat,G47gat);
xor gate_109(G341gat,G309gat,G282gat);
nand gate_110(G342gat,G319gat,G60gat);
xor gate_111(G343gat,G309gat,G285gat);
nand gate_112(G344gat,G319gat,G73gat);
nand gate_113(G345gat,G319gat,G86gat);
nand gate_114(G346gat,G319gat,G99gat);
nand gate_115(G347gat,G319gat,G112gat);
nand gate_116(G348gat,G330gat,G300gat);
nand gate_117(G349gat,G331gat,G301gat);
nand gate_118(G350gat,G332gat,G302gat);
nand gate_119(G351gat,G333gat,G303gat);
nand gate_120(G352gat,G335gat,G304gat);
nand gate_121(G353gat,G337gat,G305gat);
nand gate_122(G354gat,G339gat,G306gat);
nand gate_123(G355gat,G341gat,G307gat);
nand gate_124(G356gat,G343gat,G308gat);
and gate_125(G357gat,G348gat,G349gat,G350gat,G351gat,G352gat,G353gat,G354gat,G355gat,G356gat);
not gate_126(G360gat,G357gat);
not gate_127(G370gat,G357gat);
nand gate_128(G371gat,G14gat,G360gat);
nand gate_129(G372gat,G360gat,G27gat);
nand gate_130(G373gat,G360gat,G40gat);
nand gate_131(G374gat,G360gat,G53gat);
nand gate_132(G375gat,G360gat,G66gat);
nand gate_133(G376gat,G360gat,G79gat);
nand gate_134(G377gat,G360gat,G92gat);
nand gate_135(G378gat,G360gat,G105gat);
nand gate_136(G379gat,G360gat,G115gat);
nand gate_137(G380gat,G4gat,G242gat,G334gat,G371gat);
nand gate_138(G381gat,G246gat,G336gat,G372gat,G17gat);
nand gate_139(G386gat,G250gat,G338gat,G373gat,G30gat);
nand gate_140(G393gat,G254gat,G340gat,G374gat,G43gat);
nand gate_141(G399gat,G255gat,G342gat,G375gat,G56gat);
nand gate_142(G404gat,G256gat,G344gat,G376gat,G69gat);
nand gate_143(G407gat,G257gat,G345gat,G377gat,G82gat);
nand gate_144(G411gat,G258gat,G346gat,G378gat,G95gat);
nand gate_145(G414gat,G259gat,G347gat,G379gat,G108gat);
not gate_146(G415gat,G380gat);
and gate_147(G416gat,G381gat,G386gat,G393gat,G399gat,G404gat,G407gat,G411gat,G414gat);
not gate_148(G417gat,G393gat);
not gate_149(G418gat,G404gat);
not gate_150(G419gat,G407gat);
not gate_151(G420gat,G411gat);
nor gate_152(G421gat,G415gat,G416gat);
nand gate_153(G422gat,G386gat,G417gat);
nand gate_154(G425gat,G386gat,G393gat,G418gat,G399gat);
nand gate_155(G428gat,G399gat,G393gat,G419gat);
nand gate_156(G429gat,G386gat,G393gat,G407gat,G420gat);
nand gate_157(G430gat,G381gat,G386gat,G422gat,G399gat);
nand gate_158(G431gat,G381gat,G386gat,G425gat,G428gat);
nand gate_159(G432gat,G381gat,G422gat,G425gat,G429gat);
endmodule
