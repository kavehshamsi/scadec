// Verilog File 
module c5315 (G1,G4,G11,G14,G17,G20,G23,G24,G25,
G26,G27,G31,G34,G37,G40,G43,G46,G49,G52,
G53,G54,G61,G64,G67,G70,G73,G76,G79,G80,
G81,G82,G83,G86,G87,G88,G91,G94,G97,G100,
G103,G106,G109,G112,G113,G114,G115,G116,G117,G118,
G119,G120,G121,G122,G123,G126,G127,G128,G129,G130,
G131,G132,G135,G136,G137,G140,G141,G145,G146,G149,
G152,G155,G158,G161,G164,G167,G170,G173,G176,G179,
G182,G185,G188,G191,G194,G197,G200,G203,G206,G209,
G210,G217,G218,G225,G226,G233,G234,G241,G242,G245,
G248,G251,G254,G257,G264,G265,G272,G273,G280,G281,
G288,G289,G292,G293,G299,G302,G307,G308,G315,G316,
G323,G324,G331,G332,G335,G338,G341,G348,G351,G358,
G361,G366,G369,G372,G373,G374,G386,G389,G400,G411,
G422,G435,G446,G457,G468,G479,G490,G503,G514,G523,
G534,G545,G549,G552,G556,G559,G562,G1497,G1689,G1690,
G1691,G1694,G2174,G2358,G2824,G3173,G3546,G3548,G3550,G3552,
G3717,G3724,G4087,G4088,G4089,G4090,G4091,G4092,G4115,G144,
G298,G973,G594,G599,G600,G601,G602,G603,G604,G611,
G612,G810,G848,G849,G850,G851,G634,G815,G845,G847,
G926,G923,G921,G892,G887,G606,G656,G809,G993,G978,
G949,G939,G889,G593,G636,G704,G717,G820,G639,G673,
G707,G715,G598,G610,G588,G615,G626,G632,G1002,G1004,
G591,G618,G621,G629,G822,G838,G861,G623,G722,G832,
G834,G836,G859,G871,G873,G875,G877,G998,G1000,G575,
G585,G661,G693,G747,G752,G757,G762,G787,G792,G797,
G802,G642,G664,G667,G670,G676,G696,G699,G702,G818,
G813,G824,G826,G828,G830,G854,G863,G865,G867,G869,
G712,G727,G732,G737,G742,G772,G777,G782,G645,G648,
G651,G654,G679,G682,G685,G688,G843,G882,G767,G807,
G658,G690);

input G1,G4,G11,G14,G17,G20,G23,G24,G25,
G26,G27,G31,G34,G37,G40,G43,G46,G49,G52,
G53,G54,G61,G64,G67,G70,G73,G76,G79,G80,
G81,G82,G83,G86,G87,G88,G91,G94,G97,G100,
G103,G106,G109,G112,G113,G114,G115,G116,G117,G118,
G119,G120,G121,G122,G123,G126,G127,G128,G129,G130,
G131,G132,G135,G136,G137,G140,G141,G145,G146,G149,
G152,G155,G158,G161,G164,G167,G170,G173,G176,G179,
G182,G185,G188,G191,G194,G197,G200,G203,G206,G209,
G210,G217,G218,G225,G226,G233,G234,G241,G242,G245,
G248,G251,G254,G257,G264,G265,G272,G273,G280,G281,
G288,G289,G292,G293,G299,G302,G307,G308,G315,G316,
G323,G324,G331,G332,G335,G338,G341,G348,G351,G358,
G361,G366,G369,G372,G373,G374,G386,G389,G400,G411,
G422,G435,G446,G457,G468,G479,G490,G503,G514,G523,
G534,G545,G549,G552,G556,G559,G562,G1497,G1689,G1690,
G1691,G1694,G2174,G2358,G2824,G3173,G3546,G3548,G3550,G3552,
G3717,G3724,G4087,G4088,G4089,G4090,G4091,G4092,G4115;

output G144,G298,G973,G594,G599,G600,G601,G602,G603,
G604,G611,G612,G810,G848,G849,G850,G851,G634,G815,
G845,G847,G926,G923,G921,G892,G887,G606,G656,G809,
G993,G978,G949,G939,G889,G593,G636,G704,G717,G820,
G639,G673,G707,G715,G598,G610,G588,G615,G626,G632,
G1002,G1004,G591,G618,G621,G629,G822,G838,G861,G623,
G722,G832,G834,G836,G859,G871,G873,G875,G877,G998,
G1000,G575,G585,G661,G693,G747,G752,G757,G762,G787,
G792,G797,G802,G642,G664,G667,G670,G676,G696,G699,
G702,G818,G813,G824,G826,G828,G830,G854,G863,G865,
G867,G869,G712,G727,G732,G737,G742,G772,G777,G782,
G645,G648,G651,G654,G679,G682,G685,G688,G843,G882,
G767,G807,G658,G690;

wire G4114,G2825,G3547,G3549,G3551,G3553,G633,G814,G816,
G844,G846,G852,G1502,G1528,G1552,G1609,G1633,G1697,G1698,
G1701,G2179,G2203,G2226,G2281,G2304,G2361,G2370,G2382,G2393,
G2405,G2418,G2442,G2476,G2500,G2533,G2537,G2541,G2545,G2549,
G2553,G2557,G2561,G2627,G2631,G2635,G2639,G2643,G2647,G2651,
G2655,G2721,G2734,G2816,G2822,G2826,G2828,G2882,G2886,G2890,
G2894,G2898,G2902,G2948,G2952,G2956,G2960,G2964,G2968,G3024,
G3028,G3032,G3036,G3040,G3044,G3048,G3052,G3092,G3105,G3175,
G3176,G3181,G3204,G3208,G3212,G3216,G3220,G3224,G3256,G3260,
G3264,G3268,G3272,G3276,G3302,G3314,G3354,G3358,G3362,G3366,
G3370,G3374,G3378,G3382,G3440,G3554,G3555,G3556,G3558,G3582,
G3616,G3628,G3660,G3684,G3721,G3728,G3737,G3757,G3795,G3815,
G3972,G3991,G4030,G4049,G4110,G4119,G4127,G4135,G4143,G4151,
G4159,G4167,G4175,G4183,G4188,G4276,G4284,G4292,G4300,G4308,
G4316,G4324,G4332,G4340,G4631,G4639,G4647,G4655,G4663,G4671,
G4676,G4764,G4772,G4780,G4788,G4796,G4804,G5082,G5085,G5090,
G5093,G5098,G5101,G5108,G5111,G5332,G5335,G5340,G5343,G5348,
G5351,G5356,G5359,G5369,G2979,G2999,G1580,G1586,G1592,G1598,
G1604,G1668,G1674,G1680,G1686,G2254,G2260,G2266,G2272,G2278,
G2339,G2345,G2351,G2357,G711,G721,G726,G731,G736,G741,
G746,G751,G756,G761,G766,G771,G776,G781,G786,G791,
G796,G801,G806,G3734,G842,G858,G881,G4123,G4131,G4139,
G4147,G4155,G4163,G4171,G4179,G4187,G4194,G4282,G4290,G4298,
G4306,G4314,G4322,G4330,G4338,G4346,G1526,G1540,G1564,G1606,
G1621,G1645,G1661,G1688,G4635,G4643,G4651,G4659,G4667,G4675,
G4682,G4770,G4778,G4786,G4794,G4802,G4810,G2202,G2215,G2238,
G2279,G2293,G2316,G2332,G2430,G2454,G2488,G2512,G2536,G2540,
G2544,G2548,G2552,G2556,G2560,G2564,G2566,G2572,G2578,G2584,
G2590,G2595,G2600,G2605,G2630,G2634,G2638,G2642,G2646,G2650,
G2654,G2658,G2660,G2666,G2672,G2678,G2684,G2689,G2694,G2699,
G2728,G2741,G2748,G2750,G2752,G2754,G2756,G2758,G2760,G2762,
G2764,G2766,G2827,G2838,G2847,G2885,G2889,G2893,G2897,G2901,
G2905,G2906,G2909,G2913,G2918,G2922,G2927,G2951,G2955,G2959,
G2963,G2967,G2971,G2973,G2980,G2982,G2988,G2994,G3001,G3006,
G3027,G3031,G3035,G3039,G3043,G3047,G3051,G3055,G3056,G3060,
G3064,G3068,G3073,G3078,G3083,G3088,G3099,G3112,G3119,G3121,
G3123,G3125,G3126,G3128,G3130,G3132,G3134,G3136,G3187,G3193,
G3196,G3199,G3202,G3207,G3211,G3215,G3219,G3223,G3227,G3228,
G3232,G3234,G3238,G3243,G3247,G3249,G3253,G3259,G3263,G3267,
G3271,G3275,G3279,G3280,G3283,G3287,G3292,G3295,G3299,G3305,
G3306,G3310,G3317,G3318,G3322,G3326,G3333,G3357,G3361,G3365,
G3369,G3373,G3377,G3381,G3385,G3386,G3390,G3394,G3398,G3403,
G3408,G3413,G3418,G5088,G5089,G5096,G5097,G3489,G3493,G3570,
G3594,G3622,G3632,G3637,G3640,G3643,G3646,G3672,G3696,G3745,
G3765,G3803,G3823,G5338,G5339,G5346,G5347,G5354,G5355,G3979,
G3998,G4037,G4056,G4094,G5104,G5105,G5114,G5115,G5362,G5363,
G5366,G5373,G2568,G2574,G2580,G2586,G2592,G2597,G2602,G2607,
G2662,G2668,G2674,G2680,G2686,G2691,G2696,G2701,G2907,G2910,
G2914,G2920,G2924,G2929,G2975,G2984,G2990,G2996,G3003,G3008,
G3015,G3057,G3061,G3065,G3069,G3075,G3080,G3085,G3090,G3229,
G3233,G3235,G3239,G3244,G3250,G3254,G3281,G3284,G3288,G3293,
G3296,G3300,G3327,G3334,G3387,G3391,G3395,G3399,G3405,G3410,
G3415,G3420,G3422,G3423,G3431,G3432,G3895,G3896,G3904,G3905,
G3913,G3914,G5106,G5107,G5116,G5117,G5364,G5365,G2880,G2881,
G1579,G1585,G1591,G1597,G1603,G1667,G1673,G1679,G1685,G2876,
G2877,G2253,G2259,G2265,G2271,G2277,G2338,G2344,G2350,G2356,
G2868,G2869,G710,G2872,G2873,G720,G725,G730,G735,G740,
G745,G750,G755,G760,G765,G770,G775,G780,G785,G790,
G795,G800,G805,G841,G857,G880,G1660,G2331,G2569,G2575,
G2581,G2587,G2593,G2598,G2603,G2608,G2663,G2669,G2675,G2681,
G2687,G2692,G2697,G2702,G2747,G2749,G2751,G2753,G2755,G2757,
G2759,G2761,G2763,G2765,G2857,G2908,G2911,G2915,G2925,G2930,
G2933,G2976,G2985,G2991,G2997,G3004,G3009,G3058,G3062,G3066,
G3070,G3076,G3081,G3086,G3091,G3118,G3120,G3122,G3124,G3127,
G3129,G3131,G3133,G3135,G3147,G3192,G3195,G3198,G3201,G3230,
G3236,G3240,G3245,G3251,G3255,G3282,G3285,G3289,G3297,G3301,
G3309,G3313,G3321,G3325,G3328,G3329,G3335,G3336,G3341,G3345,
G3388,G3392,G3396,G3400,G3406,G3411,G3416,G3421,G3424,G3433,
G3492,G3496,G3780,G3783,G3786,G3789,G3838,G3841,G3844,G3847,
G3897,G3906,G3915,G4011,G4014,G4017,G4020,G4023,G4069,G4072,
G4075,G4078,G4081,G5206,G5209,G5307,G5322,G5372,G5375,G5399,
G2813,G3197,G3200,G3203,G3194,G2570,G2576,G2582,G2588,G2664,
G2670,G2676,G2682,G2767,G2772,G2776,G2780,G2784,G2788,G2794,
G2798,G2802,G2912,G2916,G2936,G2977,G2986,G2992,G3059,G3063,
G3067,G3071,G3137,G3139,G3143,G3151,G3155,G3161,G3165,G3167,
G3231,G3237,G3241,G3286,G3290,G3330,G3337,G3342,G3346,G3348,
G3352,G3389,G3393,G3397,G3401,G3845,G5126,G5178,G5325,G5374,
G2810,G635,G2878,G2879,G2874,G2875,G703,G2866,G2867,G2870,
G2871,G716,G819,G1789,G2036,G2611,G2615,G2619,G2623,G2705,
G2709,G2713,G2717,G2939,G2942,G2945,G3012,G3018,G3021,G3331,
G3338,G3343,G3347,G3428,G3437,G3514,G3836,G3852,G5311,G3901,
G3910,G3934,G3938,G4652,G4783,G5137,G5212,G5213,G5260,G5263,
G5268,G5271,G5276,G5279,G5289,G5296,G5299,G5304,G5312,G5315,
G5328,G5396,G5403,G1286,G2809,G597,G1031,G637,G671,G705,
G713,G1046,G1064,G1071,G1097,G1111,G1128,G1145,G1160,G1301,
G1318,G1324,G1341,G1359,G1382,G1404,G1412,G1704,G1712,G1724,
G1742,G1749,G1775,G1806,G1823,G1829,G1837,G1958,G1966,G1978,
G1995,G2001,G2018,G2059,G2081,G2089,G2106,G3170,G3332,G3339,
G5132,G5184,G3853,G3874,G4076,G4116,G4124,G4132,G4140,G4148,
G4156,G4164,G4172,G4180,G4228,G4279,G4287,G4295,G4303,G4311,
G4319,G4327,G4335,G4343,G4348,G4464,G4628,G4636,G4644,G4660,
G4668,G4716,G4767,G4775,G4791,G4799,G4807,G4812,G5118,G5121,
G5129,G5134,G5142,G5145,G5152,G5155,G5162,G5165,G5170,G5173,
G5181,G5186,G5189,G5196,G5199,G5214,G5215,G5329,G5330,G2807,
G2808,G2811,G2812,G2814,G2626,G2622,G2618,G2614,G2720,G2716,
G2712,G2708,G3731,G4658,G1777,G2019,G4787,G3350,G3353,G5141,
G3513,G3516,G3517,G3778,G3781,G3784,G3787,G3839,G3842,G5266,
G5267,G5274,G5275,G5302,G5303,G5310,G3891,G3937,G3941,G3955,
G3958,G4009,G4012,G4015,G4018,G4067,G4070,G4073,G4079,G5239,
G5282,G5283,G5293,G5318,G5319,G5331,G5402,G5405,G595,G596,
G607,G608,G1845,G1846,G2115,G2116,G4122,G1022,G4130,G1033,
G4138,G1051,G4146,G1079,G4154,G1088,G4162,G1099,G4170,G1115,
G4178,G1133,G4186,G1151,G4234,G1276,G4283,G1287,G4291,G1305,
G4299,G1330,G4307,G1342,G4315,G1363,G4323,G1388,G4331,G1420,
G4339,G1428,G4347,G4634,G1729,G4642,G1757,G4650,G1766,G1776,
G4666,G1793,G4674,G1811,G1849,G1852,G1875,G4722,G1982,G4771,
G2007,G4779,G2020,G2040,G4795,G2065,G4803,G2097,G4811,G2119,
G2122,G5124,G5125,G3452,G5133,G5140,G3462,G5168,G5169,G5176,
G5177,G3484,G5185,G3515,G3518,G3857,G3860,G3861,G3869,G3870,
G3878,G3881,G3882,G3890,G3954,G3957,G4021,G4099,G4236,G4354,
G4406,G4470,G4552,G4679,G4687,G4695,G4703,G4711,G4724,G4818,
G4855,G4865,G4870,G4913,G4923,G4951,G5006,G5039,G5148,G5149,
G5158,G5159,G5192,G5193,G5202,G5203,G5284,G5285,G5320,G5321,
G5386,G5404,G609,G1021,G1032,G1050,G1078,G1087,G1098,G1114,
G1132,G1150,G1277,G1288,G1306,G1331,G1343,G1364,G1389,G1421,
G1429,G1728,G1756,G1765,G1778,G1792,G1810,G1983,G2008,G2021,
G2041,G2066,G2098,G3443,G3444,G3453,G3461,G3466,G3467,G3475,
G3476,G3485,G5243,G3862,G3871,G3883,G3892,G3956,G3959,G4756,
G5150,G5151,G5160,G5161,G5194,G5195,G5204,G5205,G5236,G5286,
G5379,G5389,G5425,G1023,G1034,G1052,G1080,G1089,G1100,G1116,
G1134,G1152,G4242,G1278,G1289,G1307,G1332,G1344,G1365,G1390,
G1422,G1430,G1730,G1758,G1767,G1794,G1812,G1876,G4683,G4691,
G4699,G4707,G4715,G4730,G1984,G2009,G2042,G2067,G2099,G4869,
G4927,G3445,G3454,G3463,G3468,G3477,G3486,G4103,G4412,G4558,
G4859,G4876,G4917,G4955,G5012,G5043,G5216,G5219,G5226,G5229,
G5392,G5422,G1866,G1877,G4762,G2142,G2146,G5242,G3532,G3866,
G3887,G3918,G3922,G3926,G3930,G5429,G4104,G4743,G4991,G5001,
G5292,G5295,G5383,G5393,G5394,G1439,G1440,G1441,G1847,G1168,
G1169,G1170,G2117,G1086,G1166,G1171,G1172,G1173,G1174,G1175,
G1176,G1177,G1178,G1179,G1181,G1182,G1183,G1184,G1188,G1189,
G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1437,G1442,
G1443,G1444,G1445,G1446,G1447,G1451,G1454,G1455,G1456,G1457,
G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,
G1475,G1476,G1477,G1481,G1482,G1764,G1843,G1850,G1851,G1853,
G1854,G1855,G1856,G1857,G1859,G1860,G1861,G1862,G1867,G1868,
G1869,G1870,G1871,G1872,G1873,G1874,G1878,G2113,G2120,G2121,
G2123,G2124,G2128,G2131,G2132,G2133,G2134,G2143,G2144,G2145,
G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2158,G2159,
G3449,G3458,G3472,G3481,G3497,G3501,G3505,G3509,G3531,G5428,
G3967,G4191,G4199,G4207,G4215,G4223,G4231,G4239,G4247,G4255,
G4263,G4271,G4371,G4381,G4391,G4401,G4429,G4439,G4449,G4459,
G4497,G4507,G4517,G4527,G4537,G4547,G4585,G4595,G4605,G4615,
G4719,G4727,G4735,G4751,G4759,G4835,G4845,G4893,G4903,G4961,
G4971,G4981,G5049,G5059,G5069,G5222,G5223,G5232,G5233,G5294,
G5395,G589,G616,G619,G627,G1185,G1448,G1458,G1478,G1863,
G4747,G2125,G2135,G2155,G4995,G5005,G3533,G3921,G3925,G3929,
G3933,G3943,G3946,G3949,G3952,G3966,G4107,G4196,G4204,G4212,
G4220,G4244,G4252,G4260,G4268,G4361,G4419,G4467,G4487,G4555,
G4575,G4684,G4692,G4700,G4708,G4732,G4740,G4748,G4825,G4883,
G4928,G4941,G5009,G5029,G5224,G5225,G5234,G5235,G5376,G5417,
G576,G1198,G4195,G4203,G4211,G4219,G4227,G1217,G4235,G1221,
G4243,G1224,G4251,G4259,G4267,G4275,G1453,G4405,G4463,G4541,
G4551,G1895,G4723,G1899,G4731,G1902,G4739,G4755,G1929,G4763,
G2130,G3500,G3504,G3508,G3512,G3520,G3523,G3526,G3529,G3837,
G3942,G3945,G3948,G3951,G3968,G4375,G4385,G4395,G4433,G4443,
G4453,G4501,G4511,G4521,G4531,G4619,G4589,G4599,G4609,G4839,
G4849,G4897,G4907,G4965,G4975,G4985,G5073,G5053,G5063,G5247,
G5255,G590,G617,G620,G628,G3535,G1199,G4202,G1204,G4210,
G1207,G4218,G1211,G4226,G1214,G1218,G1222,G1225,G4250,G1237,
G4258,G1242,G4266,G1247,G4274,G1252,G1462,G4690,G1882,G4698,
G1885,G4706,G1889,G4714,G1892,G1896,G1900,G1903,G4738,G1915,
G4746,G1920,G4754,G1925,G1930,G2139,G3519,G3522,G3525,G3528,
G3848,G3944,G3947,G3950,G3953,G5421,G4111,G4112,G4351,G4365,
G4409,G4423,G4471,G4472,G4477,G4491,G4559,G4560,G4565,G4579,
G4815,G4829,G4873,G4887,G4931,G4934,G4945,G5013,G5014,G5019,
G5033,G5382,G5385,G3970,G1200,G1203,G1206,G1210,G1213,G1219,
G1223,G1236,G1241,G1246,G1251,G1881,G1884,G1888,G1891,G1897,
G1901,G1914,G1919,G1924,G1931,G3521,G3524,G3527,G3530,G5251,
G5259,G4113,G4473,G4561,G5015,G5384,G5406,G5414,G1664,G2335,
G718,G855,G1205,G1208,G1212,G1215,G1220,G1231,G1238,G1243,
G1248,G1253,G1272,G1483,G1883,G1886,G1890,G1893,G1898,G1909,
G1916,G1921,G1926,G1953,G2160,G4355,G4356,G4413,G4414,G4474,
G4481,G4562,G4569,G4819,G4820,G4877,G4878,G4935,G4936,G5016,
G5023,G5244,G5252,G5409,G566,G577,G3733,G1209,G1216,G1257,
G1262,G1267,G1887,G1894,G1935,G1943,G1948,G3779,G3840,G5412,
G5420,G3964,G4357,G4415,G4821,G4879,G4937,G567,G568,G569,
G570,G578,G579,G580,G1256,G1261,G1266,G1271,G1486,G1934,
G1942,G1947,G1952,G2163,G5250,G3537,G5258,G3542,G3782,G3785,
G3788,G3790,G3843,G3846,G3849,G3960,G5413,G3963,G4010,G4068,
G4358,G4416,G4480,G4483,G4568,G4571,G4822,G4880,G4938,G5022,
G5025,G1258,G1263,G1268,G1273,G1936,G1944,G1949,G1954,G3536,
G3541,G3791,G3792,G3793,G3850,G3851,G3961,G3965,G4024,G4082,
G4482,G4570,G5024,G1666,G1670,G2337,G2341,G719,G758,G798,
G856,G3538,G3543,G3962,G4364,G4367,G4422,G4425,G4484,G4572,
G4828,G4831,G4886,G4889,G4944,G4947,G5026,G571,G572,G573,
G574,G581,G582,G583,G584,G1576,G1578,G659,G1672,G1676,
G1678,G1682,G1684,G2250,G2252,G691,G2343,G2347,G2349,G2353,
G2355,G743,G744,G748,G749,G753,G754,G759,G783,G784,
G788,G789,G793,G794,G799,G3735,G3835,G3651,G4013,G4016,
G4019,G4022,G4071,G4074,G4077,G4080,G4096,G4366,G4424,G4830,
G4888,G4946,G640,G662,G665,G668,G674,G694,G697,G700,
G817,G839,G3540,G3545,G3777,G3648,G4025,G4026,G4027,G4028,
G4083,G4084,G4085,G4086,G4368,G4426,G4490,G4493,G4578,G4581,
G4832,G4890,G4948,G5032,G5035,G811,G812,G853,G878,G4492,
G4580,G5034,G1582,G1584,G1588,G1590,G1594,G1596,G1600,G1602,
G2256,G2258,G2262,G2264,G2268,G2270,G2274,G2276,G708,G709,
G723,G724,G728,G729,G733,G734,G738,G739,G768,G769,
G773,G774,G778,G779,G4374,G4377,G4432,G4435,G4494,G4582,
G4838,G4841,G4896,G4899,G4954,G4957,G5036,G643,G646,G649,
G652,G677,G680,G683,G686,G4376,G4434,G4840,G4898,G4956,
G4378,G4436,G4500,G4503,G4588,G4591,G4842,G4900,G4958,G5042,
G5045,G4502,G4590,G5044,G4384,G4387,G4442,G4445,G4504,G4592,
G4848,G4851,G4906,G4909,G4964,G4967,G5046,G4386,G4444,G4850,
G4908,G4966,G4388,G4446,G4510,G4513,G4598,G4601,G4852,G4910,
G4968,G5052,G5055,G4512,G4600,G5054,G4394,G4397,G4452,G4455,
G4514,G4602,G4858,G4861,G4916,G4919,G4974,G4977,G5056,G4396,
G4454,G4860,G4918,G4976,G4398,G4456,G4520,G4523,G4608,G4611,
G4862,G4920,G4978,G5062,G5065,G4522,G4610,G5064,G4404,G1488,
G4462,G1493,G4868,G2165,G4926,G2170,G4524,G4612,G4984,G4987,
G5066,G1487,G1492,G2164,G2169,G4986,G1489,G1494,G2166,G2171,
G4530,G4533,G4618,G4543,G4988,G5072,G4997,G4532,G4542,G4996,
G1513,G1514,G1515,G1516,G4994,G2184,G2190,G2191,G2192,G2193,
G4534,G4544,G4998,G2183,G4620,G5074,G4540,G1507,G4550,G1510,
G2185,G5004,G2187,G1506,G1509,G4626,G2186,G2195,G5080,G1508,
G1511,G2188,G1512,G1518,G2189,G1517,G2194,G4623,G5077,G1519,
G4627,G2196,G5081,G1520,G2197,G1521,G2198,G840,G879,G1524,
G2201,G3649,G3652,G3657,G3658,G3636,G3639,G3642,G3645,G3653,
G3654,G3655,G3656,G763,G764,G803,G804,G1657,G1659,G2328,
G2330,G1662,G2333,G657,G689;
buf gate_0(G144,G141);
buf gate_1(G298,G293);
and gate_2(G4114,G135,G4115);
not gate_3(G2825,G2824);
buf gate_4(G973,G3173);
not gate_5(G3547,G3546);
not gate_6(G3549,G3548);
not gate_7(G3551,G3550);
not gate_8(G3553,G3552);
not gate_9(G594,G545);
not gate_10(G599,G348);
not gate_11(G600,G366);
and gate_12(G601,G552,G562);
not gate_13(G602,G549);
not gate_14(G603,G545);
not gate_15(G604,G545);
not gate_16(G611,G338);
not gate_17(G612,G358);
nand gate_18(G633,G373,G1);
and gate_19(G810,G141,G145);
not gate_20(G814,G3173);
not gate_21(G816,G4114);
and gate_22(G844,G2825,G27);
and gate_23(G846,G386,G556);
not gate_24(G848,G245);
not gate_25(G849,G552);
not gate_26(G850,G562);
not gate_27(G851,G559);
and gate_28(G852,G386,G559,G556,G552);
not gate_29(G1502,G1497);
buf gate_30(G1528,G1689);
buf gate_31(G1552,G1690);
buf gate_32(G1609,G1689);
buf gate_33(G1633,G1690);
buf gate_34(G1697,G137);
buf gate_35(G1698,G137);
buf gate_36(G1701,G141);
not gate_37(G2179,G2174);
buf gate_38(G2203,G1691);
buf gate_39(G2226,G1694);
buf gate_40(G2281,G1691);
buf gate_41(G2304,G1694);
buf gate_42(G2361,G254);
buf gate_43(G2370,G251);
buf gate_44(G2382,G251);
buf gate_45(G2393,G248);
buf gate_46(G2405,G248);
buf gate_47(G2418,G4088);
buf gate_48(G2442,G4087);
buf gate_49(G2476,G4089);
buf gate_50(G2500,G4090);
buf gate_51(G2533,G210);
buf gate_52(G2537,G210);
buf gate_53(G2541,G218);
buf gate_54(G2545,G218);
buf gate_55(G2549,G226);
buf gate_56(G2553,G226);
buf gate_57(G2557,G234);
buf gate_58(G2561,G234);
buf gate_59(G2627,G257);
buf gate_60(G2631,G257);
buf gate_61(G2635,G265);
buf gate_62(G2639,G265);
buf gate_63(G2643,G273);
buf gate_64(G2647,G273);
buf gate_65(G2651,G281);
buf gate_66(G2655,G281);
buf gate_67(G2721,G335);
buf gate_68(G2734,G335);
buf gate_69(G2816,G206);
and gate_70(G2822,G27,G31);
buf gate_71(G2826,G1);
buf gate_72(G2828,G2358);
buf gate_73(G2882,G293);
buf gate_74(G2886,G302);
buf gate_75(G2890,G308);
buf gate_76(G2894,G308);
buf gate_77(G2898,G316);
buf gate_78(G2902,G316);
buf gate_79(G2948,G324);
buf gate_80(G2952,G324);
buf gate_81(G2956,G341);
buf gate_82(G2960,G341);
buf gate_83(G2964,G351);
buf gate_84(G2968,G351);
buf gate_85(G3024,G257);
buf gate_86(G3028,G257);
buf gate_87(G3032,G265);
buf gate_88(G3036,G265);
buf gate_89(G3040,G273);
buf gate_90(G3044,G273);
buf gate_91(G3048,G281);
buf gate_92(G3052,G281);
buf gate_93(G3092,G332);
buf gate_94(G3105,G332);
buf gate_95(G3175,G549);
and gate_96(G3176,G31,G27);
not gate_97(G3181,G2358);
buf gate_98(G3204,G324);
buf gate_99(G3208,G324);
buf gate_100(G3212,G341);
buf gate_101(G3216,G341);
buf gate_102(G3220,G351);
buf gate_103(G3224,G351);
buf gate_104(G3256,G293);
buf gate_105(G3260,G302);
buf gate_106(G3264,G308);
buf gate_107(G3268,G308);
buf gate_108(G3272,G316);
buf gate_109(G3276,G316);
buf gate_110(G3302,G361);
buf gate_111(G3314,G361);
buf gate_112(G3354,G210);
buf gate_113(G3358,G210);
buf gate_114(G3362,G218);
buf gate_115(G3366,G218);
buf gate_116(G3370,G226);
buf gate_117(G3374,G226);
buf gate_118(G3378,G234);
buf gate_119(G3382,G234);
not gate_120(G3440,G324);
buf gate_121(G3554,G242);
buf gate_122(G3555,G242);
buf gate_123(G3556,G254);
buf gate_124(G3558,G4088);
buf gate_125(G3582,G4087);
buf gate_126(G3616,G4092);
buf gate_127(G3628,G4091);
buf gate_128(G3660,G4089);
buf gate_129(G3684,G4090);
not gate_130(G3721,G3717);
not gate_131(G3728,G3724);
buf gate_132(G3737,G4091);
buf gate_133(G3757,G4092);
buf gate_134(G3795,G4091);
buf gate_135(G3815,G4092);
buf gate_136(G3972,G4091);
buf gate_137(G3991,G4092);
buf gate_138(G4030,G4091);
buf gate_139(G4049,G4092);
buf gate_140(G4110,G299);
buf gate_141(G4119,G446);
buf gate_142(G4127,G457);
buf gate_143(G4135,G468);
buf gate_144(G4143,G422);
buf gate_145(G4151,G435);
buf gate_146(G4159,G389);
buf gate_147(G4167,G400);
buf gate_148(G4175,G411);
buf gate_149(G4183,G374);
buf gate_150(G4188,G4);
buf gate_151(G4276,G446);
buf gate_152(G4284,G457);
buf gate_153(G4292,G468);
buf gate_154(G4300,G435);
buf gate_155(G4308,G389);
buf gate_156(G4316,G400);
buf gate_157(G4324,G411);
buf gate_158(G4332,G422);
buf gate_159(G4340,G374);
buf gate_160(G4631,G479);
buf gate_161(G4639,G490);
buf gate_162(G4647,G503);
buf gate_163(G4655,G514);
buf gate_164(G4663,G523);
buf gate_165(G4671,G534);
buf gate_166(G4676,G54);
buf gate_167(G4764,G479);
buf gate_168(G4772,G503);
buf gate_169(G4780,G514);
buf gate_170(G4788,G523);
buf gate_171(G4796,G534);
buf gate_172(G4804,G490);
buf gate_173(G5082,G361);
buf gate_174(G5085,G369);
buf gate_175(G5090,G341);
buf gate_176(G5093,G351);
buf gate_177(G5098,G308);
buf gate_178(G5101,G316);
buf gate_179(G5108,G293);
buf gate_180(G5111,G302);
buf gate_181(G5332,G281);
buf gate_182(G5335,G289);
buf gate_183(G5340,G265);
buf gate_184(G5343,G273);
buf gate_185(G5348,G234);
buf gate_186(G5351,G257);
buf gate_187(G5356,G218);
buf gate_188(G5359,G226);
buf gate_189(G5369,G210);
not gate_190(G634,G633);
and gate_191(G815,G136,G814);
not gate_192(G845,G844);
not gate_193(G847,G846);
buf gate_194(G926,G1697);
buf gate_195(G923,G1701);
buf gate_196(G921,G2826);
and gate_197(G2979,G3553,G514);
or gate_198(G2999,G3547,G514);
buf gate_199(G892,G3175);
buf gate_200(G887,G4110);
not gate_201(G606,G3175);
and gate_202(G1580,G170,G1528,G1552);
and gate_203(G1586,G173,G1528,G1552);
and gate_204(G1592,G167,G1528,G1552);
and gate_205(G1598,G164,G1528,G1552);
and gate_206(G1604,G161,G1528,G1552);
nand gate_207(G656,G2822,G140);
and gate_208(G1668,G185,G1609,G1633);
and gate_209(G1674,G158,G1609,G1633);
and gate_210(G1680,G152,G1609,G1633);
and gate_211(G1686,G146,G1609,G1633);
and gate_212(G2254,G170,G2203,G2226);
and gate_213(G2260,G173,G2203,G2226);
and gate_214(G2266,G167,G2203,G2226);
and gate_215(G2272,G164,G2203,G2226);
and gate_216(G2278,G161,G2203,G2226);
and gate_217(G2339,G185,G2281,G2304);
and gate_218(G2345,G158,G2281,G2304);
and gate_219(G2351,G152,G2281,G2304);
and gate_220(G2357,G146,G2281,G2304);
and gate_221(G711,G106,G3660,G3684);
and gate_222(G721,G61,G2418,G2442);
and gate_223(G726,G106,G3558,G3582);
and gate_224(G731,G49,G3558,G3582);
and gate_225(G736,G103,G3558,G3582);
and gate_226(G741,G40,G3558,G3582);
and gate_227(G746,G37,G3558,G3582);
and gate_228(G751,G20,G2418,G2442);
and gate_229(G756,G17,G2418,G2442);
and gate_230(G761,G70,G2418,G2442);
and gate_231(G766,G64,G2418,G2442);
and gate_232(G771,G49,G3660,G3684);
and gate_233(G776,G103,G3660,G3684);
and gate_234(G781,G40,G3660,G3684);
and gate_235(G786,G37,G3660,G3684);
and gate_236(G791,G20,G2476,G2500);
and gate_237(G796,G17,G2476,G2500);
and gate_238(G801,G70,G2476,G2500);
and gate_239(G806,G64,G2476,G2500);
not gate_240(G809,G2822);
and gate_241(G3734,G123,G3728,G3717);
and gate_242(G842,G3795,G3815);
and gate_243(G858,G61,G2476,G2500);
and gate_244(G881,G3737,G3757);
not gate_245(G4123,G4119);
not gate_246(G4131,G4127);
not gate_247(G4139,G4135);
not gate_248(G4147,G4143);
not gate_249(G4155,G4151);
not gate_250(G4163,G4159);
not gate_251(G4171,G4167);
not gate_252(G4179,G4175);
not gate_253(G4187,G4183);
not gate_254(G4194,G4188);
not gate_255(G4282,G4276);
not gate_256(G4290,G4284);
not gate_257(G4298,G4292);
not gate_258(G4306,G4300);
not gate_259(G4314,G4308);
not gate_260(G4322,G4316);
not gate_261(G4330,G4324);
not gate_262(G4338,G4332);
not gate_263(G4346,G4340);
buf gate_264(G1526,G1697);
not gate_265(G1540,G1528);
not gate_266(G1564,G1552);
buf gate_267(G1606,G1697);
not gate_268(G1621,G1609);
not gate_269(G1645,G1633);
and gate_270(G1661,G179,G1609,G1633);
buf gate_271(G1688,G2826);
not gate_272(G4635,G4631);
not gate_273(G4643,G4639);
not gate_274(G4651,G4647);
not gate_275(G4659,G4655);
not gate_276(G4667,G4663);
not gate_277(G4675,G4671);
not gate_278(G4682,G4676);
not gate_279(G4770,G4764);
not gate_280(G4778,G4772);
not gate_281(G4786,G4780);
not gate_282(G4794,G4788);
not gate_283(G4802,G4796);
not gate_284(G4810,G4804);
buf gate_285(G2202,G1698);
not gate_286(G2215,G2203);
not gate_287(G2238,G2226);
buf gate_288(G2279,G1698);
not gate_289(G2293,G2281);
not gate_290(G2316,G2304);
and gate_291(G2332,G179,G2281,G2304);
not gate_292(G2430,G2418);
not gate_293(G2454,G2442);
not gate_294(G2488,G2476);
not gate_295(G2512,G2500);
not gate_296(G2536,G2533);
not gate_297(G2540,G2537);
not gate_298(G2544,G2541);
not gate_299(G2548,G2545);
not gate_300(G2552,G2549);
not gate_301(G2556,G2553);
not gate_302(G2560,G2557);
not gate_303(G2564,G2561);
and gate_304(G2566,G3553,G457,G2537);
and gate_305(G2572,G3553,G468,G2545);
and gate_306(G2578,G3553,G422,G2553);
and gate_307(G2584,G3553,G435,G2561);
and gate_308(G2590,G3547,G2533);
and gate_309(G2595,G3547,G2541);
and gate_310(G2600,G3547,G2549);
and gate_311(G2605,G3547,G2557);
not gate_312(G2630,G2627);
not gate_313(G2634,G2631);
not gate_314(G2638,G2635);
not gate_315(G2642,G2639);
not gate_316(G2646,G2643);
not gate_317(G2650,G2647);
not gate_318(G2654,G2651);
not gate_319(G2658,G2655);
and gate_320(G2660,G3553,G389,G2631);
and gate_321(G2666,G3553,G400,G2639);
and gate_322(G2672,G3553,G411,G2647);
and gate_323(G2678,G3553,G374,G2655);
and gate_324(G2684,G3547,G2627);
and gate_325(G2689,G3547,G2635);
and gate_326(G2694,G3547,G2643);
and gate_327(G2699,G3547,G2651);
not gate_328(G2728,G2721);
not gate_329(G2741,G2734);
and gate_330(G2748,G292,G2721);
and gate_331(G2750,G288,G2721);
and gate_332(G2752,G280,G2721);
and gate_333(G2754,G272,G2721);
and gate_334(G2756,G264,G2721);
and gate_335(G2758,G241,G2734);
and gate_336(G2760,G233,G2734);
and gate_337(G2762,G225,G2734);
and gate_338(G2764,G217,G2734);
and gate_339(G2766,G209,G2734);
buf gate_340(G2827,G1701);
not gate_341(G2838,G2828);
not gate_342(G2847,G2822);
not gate_343(G2885,G2882);
not gate_344(G2889,G2886);
not gate_345(G2893,G2890);
not gate_346(G2897,G2894);
not gate_347(G2901,G2898);
not gate_348(G2905,G2902);
and gate_349(G2906,G2393,G2886);
and gate_350(G2909,G2393,G479,G2894);
and gate_351(G2913,G2393,G490,G2902);
and gate_352(G2918,G3554,G2882);
and gate_353(G2922,G3554,G2890);
and gate_354(G2927,G3554,G2898);
not gate_355(G2951,G2948);
not gate_356(G2955,G2952);
not gate_357(G2959,G2956);
not gate_358(G2963,G2960);
not gate_359(G2967,G2964);
not gate_360(G2971,G2968);
and gate_361(G2973,G3553,G503,G2952);
not gate_362(G2980,G2979);
and gate_363(G2982,G3553,G523,G2960);
and gate_364(G2988,G3553,G534,G2968);
and gate_365(G2994,G3547,G2948);
and gate_366(G3001,G3547,G2956);
and gate_367(G3006,G3547,G2964);
not gate_368(G3027,G3024);
not gate_369(G3031,G3028);
not gate_370(G3035,G3032);
not gate_371(G3039,G3036);
not gate_372(G3043,G3040);
not gate_373(G3047,G3044);
not gate_374(G3051,G3048);
not gate_375(G3055,G3052);
and gate_376(G3056,G2393,G389,G3028);
and gate_377(G3060,G2393,G400,G3036);
and gate_378(G3064,G2393,G411,G3044);
and gate_379(G3068,G2393,G374,G3052);
and gate_380(G3073,G3554,G3024);
and gate_381(G3078,G3554,G3032);
and gate_382(G3083,G3554,G3040);
and gate_383(G3088,G3554,G3048);
not gate_384(G3099,G3092);
not gate_385(G3112,G3105);
and gate_386(G3119,G372,G3092);
and gate_387(G3121,G366,G3092);
and gate_388(G3123,G358,G3092);
and gate_389(G3125,G348,G3092);
and gate_390(G3126,G338,G3092);
and gate_391(G3128,G331,G3105);
and gate_392(G3130,G323,G3105);
and gate_393(G3132,G315,G3105);
and gate_394(G3134,G307,G3105);
and gate_395(G3136,G299,G3105);
not gate_396(G3187,G3181);
and gate_397(G3193,G83,G3181);
and gate_398(G3196,G86,G3181);
and gate_399(G3199,G88,G3181);
and gate_400(G3202,G88,G3181);
not gate_401(G3207,G3204);
not gate_402(G3211,G3208);
not gate_403(G3215,G3212);
not gate_404(G3219,G3216);
not gate_405(G3223,G3220);
not gate_406(G3227,G3224);
and gate_407(G3228,G2405,G503,G3208);
and gate_408(G3232,G2405,G514);
and gate_409(G3234,G2405,G523,G3216);
and gate_410(G3238,G2405,G534,G3224);
and gate_411(G3243,G3555,G3204);
or gate_412(G3247,G3555,G514);
and gate_413(G3249,G3555,G3212);
and gate_414(G3253,G3555,G3220);
not gate_415(G3259,G3256);
not gate_416(G3263,G3260);
not gate_417(G3267,G3264);
not gate_418(G3271,G3268);
not gate_419(G3275,G3272);
not gate_420(G3279,G3276);
and gate_421(G3280,G2405,G3260);
and gate_422(G3283,G2405,G479,G3268);
and gate_423(G3287,G2405,G490,G3276);
and gate_424(G3292,G3555,G3256);
and gate_425(G3295,G3555,G3264);
and gate_426(G3299,G3555,G3272);
not gate_427(G3305,G3302);
buf gate_428(G3306,G2816);
buf gate_429(G3310,G2816);
not gate_430(G3317,G3314);
buf gate_431(G3318,G2816);
buf gate_432(G3322,G2816);
and gate_433(G3326,G2405,G3302);
and gate_434(G3333,G2405,G3314);
not gate_435(G3357,G3354);
not gate_436(G3361,G3358);
not gate_437(G3365,G3362);
not gate_438(G3369,G3366);
not gate_439(G3373,G3370);
not gate_440(G3377,G3374);
not gate_441(G3381,G3378);
not gate_442(G3385,G3382);
and gate_443(G3386,G2393,G457,G3358);
and gate_444(G3390,G2393,G468,G3366);
and gate_445(G3394,G2393,G422,G3374);
and gate_446(G3398,G2393,G435,G3382);
and gate_447(G3403,G3554,G3354);
and gate_448(G3408,G3554,G3362);
and gate_449(G3413,G3554,G3370);
and gate_450(G3418,G3554,G3378);
not gate_451(G5088,G5082);
not gate_452(G5089,G5085);
not gate_453(G5096,G5090);
not gate_454(G5097,G5093);
buf gate_455(G3489,G3440);
buf gate_456(G3493,G3440);
not gate_457(G3570,G3558);
not gate_458(G3594,G3582);
not gate_459(G3622,G3616);
not gate_460(G3632,G3628);
and gate_461(G3637,G97,G3616);
and gate_462(G3640,G94,G3616);
and gate_463(G3643,G97,G3616);
and gate_464(G3646,G94,G3616);
not gate_465(G3672,G3660);
not gate_466(G3696,G3684);
not gate_467(G3745,G3737);
not gate_468(G3765,G3757);
not gate_469(G3803,G3795);
not gate_470(G3823,G3815);
not gate_471(G5338,G5332);
not gate_472(G5339,G5335);
not gate_473(G5346,G5340);
not gate_474(G5347,G5343);
not gate_475(G5354,G5348);
not gate_476(G5355,G5351);
not gate_477(G3979,G3972);
not gate_478(G3998,G3991);
not gate_479(G4037,G4030);
not gate_480(G4056,G4049);
buf gate_481(G4094,G4110);
not gate_482(G5104,G5098);
not gate_483(G5105,G5101);
not gate_484(G5114,G5108);
not gate_485(G5115,G5111);
not gate_486(G5362,G5356);
not gate_487(G5363,G5359);
buf gate_488(G5366,G2816);
not gate_489(G5373,G5369);
buf gate_490(G993,G1688);
buf gate_491(G978,G1688);
buf gate_492(G949,G1688);
buf gate_493(G939,G1688);
and gate_494(G2568,G457,G3551,G2540);
and gate_495(G2574,G468,G3551,G2548);
and gate_496(G2580,G422,G3551,G2556);
and gate_497(G2586,G435,G3551,G2564);
and gate_498(G2592,G3549,G2536);
and gate_499(G2597,G3549,G2544);
and gate_500(G2602,G3549,G2552);
and gate_501(G2607,G3549,G2560);
and gate_502(G2662,G389,G3551,G2634);
and gate_503(G2668,G400,G3551,G2642);
and gate_504(G2674,G411,G3551,G2650);
and gate_505(G2680,G374,G3551,G2658);
and gate_506(G2686,G3549,G2630);
and gate_507(G2691,G3549,G2638);
and gate_508(G2696,G3549,G2646);
and gate_509(G2701,G3549,G2654);
and gate_510(G2907,G2370,G2889);
and gate_511(G2910,G479,G2370,G2897);
and gate_512(G2914,G490,G2370,G2905);
and gate_513(G2920,G3556,G2885);
and gate_514(G2924,G3556,G2893);
and gate_515(G2929,G3556,G2901);
and gate_516(G2975,G503,G3551,G2955);
and gate_517(G2984,G523,G3551,G2963);
and gate_518(G2990,G534,G3551,G2971);
and gate_519(G2996,G3549,G2951);
and gate_520(G3003,G3549,G2959);
and gate_521(G3008,G3549,G2967);
and gate_522(G3015,G2980,G2999);
and gate_523(G3057,G389,G2370,G3031);
and gate_524(G3061,G400,G2370,G3039);
and gate_525(G3065,G411,G2370,G3047);
and gate_526(G3069,G374,G2370,G3055);
and gate_527(G3075,G3556,G3027);
and gate_528(G3080,G3556,G3035);
and gate_529(G3085,G3556,G3043);
and gate_530(G3090,G3556,G3051);
and gate_531(G3229,G503,G2382,G3211);
not gate_532(G3233,G3232);
and gate_533(G3235,G523,G2382,G3219);
and gate_534(G3239,G534,G2382,G3227);
and gate_535(G3244,G2361,G3207);
and gate_536(G3250,G2361,G3215);
and gate_537(G3254,G2361,G3223);
and gate_538(G3281,G2382,G3263);
and gate_539(G3284,G479,G2382,G3271);
and gate_540(G3288,G490,G2382,G3279);
and gate_541(G3293,G2361,G3259);
and gate_542(G3296,G2361,G3267);
and gate_543(G3300,G2361,G3275);
and gate_544(G3327,G2382,G3305);
and gate_545(G3334,G2382,G3317);
and gate_546(G3387,G457,G2370,G3361);
and gate_547(G3391,G468,G2370,G3369);
and gate_548(G3395,G422,G2370,G3377);
and gate_549(G3399,G435,G2370,G3385);
and gate_550(G3405,G3556,G3357);
and gate_551(G3410,G3556,G3365);
and gate_552(G3415,G3556,G3373);
and gate_553(G3420,G3556,G3381);
nand gate_554(G3422,G5085,G5088);
nand gate_555(G3423,G5082,G5089);
nand gate_556(G3431,G5093,G5096);
nand gate_557(G3432,G5090,G5097);
nand gate_558(G3895,G5335,G5338);
nand gate_559(G3896,G5332,G5339);
nand gate_560(G3904,G5343,G5346);
nand gate_561(G3905,G5340,G5347);
nand gate_562(G3913,G5351,G5354);
nand gate_563(G3914,G5348,G5355);
buf gate_564(G889,G4094);
nand gate_565(G5106,G5101,G5104);
nand gate_566(G5107,G5098,G5105);
nand gate_567(G5116,G5111,G5114);
nand gate_568(G5117,G5108,G5115);
nand gate_569(G5364,G5359,G5362);
nand gate_570(G5365,G5356,G5363);
not gate_571(G593,G4094);
and gate_572(G2880,G2838,G2847);
and gate_573(G2881,G2828,G2847);
and gate_574(G1579,G200,G1540,G1552);
and gate_575(G1585,G203,G1540,G1552);
and gate_576(G1591,G197,G1540,G1552);
and gate_577(G1597,G194,G1540,G1552);
and gate_578(G1603,G191,G1540,G1552);
and gate_579(G1667,G182,G1621,G1633);
and gate_580(G1673,G188,G1621,G1633);
and gate_581(G1679,G155,G1621,G1633);
and gate_582(G1685,G149,G1621,G1633);
and gate_583(G2876,G2838,G2847);
and gate_584(G2877,G2828,G2847);
and gate_585(G2253,G200,G2215,G2226);
and gate_586(G2259,G203,G2215,G2226);
and gate_587(G2265,G197,G2215,G2226);
and gate_588(G2271,G194,G2215,G2226);
and gate_589(G2277,G191,G2215,G2226);
and gate_590(G2338,G182,G2293,G2304);
and gate_591(G2344,G188,G2293,G2304);
and gate_592(G2350,G155,G2293,G2304);
and gate_593(G2356,G149,G2293,G2304);
and gate_594(G2868,G2838,G2847);
and gate_595(G2869,G2828,G2847);
and gate_596(G710,G109,G3672,G3684);
and gate_597(G2872,G2838,G2847);
and gate_598(G2873,G2828,G2847);
and gate_599(G720,G11,G2430,G2442);
and gate_600(G725,G109,G3570,G3582);
and gate_601(G730,G46,G3570,G3582);
and gate_602(G735,G100,G3570,G3582);
and gate_603(G740,G91,G3570,G3582);
and gate_604(G745,G43,G3570,G3582);
and gate_605(G750,G76,G2430,G2442);
and gate_606(G755,G73,G2430,G2442);
and gate_607(G760,G67,G2430,G2442);
and gate_608(G765,G14,G2430,G2442);
and gate_609(G770,G46,G3672,G3684);
and gate_610(G775,G100,G3672,G3684);
and gate_611(G780,G91,G3672,G3684);
and gate_612(G785,G43,G3672,G3684);
and gate_613(G790,G76,G2488,G2500);
and gate_614(G795,G73,G2488,G2500);
and gate_615(G800,G67,G2488,G2500);
and gate_616(G805,G14,G2488,G2500);
and gate_617(G841,G120,G3803,G3815);
and gate_618(G857,G11,G2488,G2500);
and gate_619(G880,G118,G3745,G3757);
and gate_620(G1660,G176,G1621,G1633);
and gate_621(G2331,G176,G2293,G2304);
or gate_622(G2569,G2566,G2568);
or gate_623(G2575,G2572,G2574);
or gate_624(G2581,G2578,G2580);
or gate_625(G2587,G2584,G2586);
or gate_626(G2593,G2590,G2592,G457);
or gate_627(G2598,G2595,G2597,G468);
or gate_628(G2603,G2600,G2602,G422);
or gate_629(G2608,G2605,G2607,G435);
or gate_630(G2663,G2660,G2662);
or gate_631(G2669,G2666,G2668);
or gate_632(G2675,G2672,G2674);
or gate_633(G2681,G2678,G2680);
or gate_634(G2687,G2684,G2686,G389);
or gate_635(G2692,G2689,G2691,G400);
or gate_636(G2697,G2694,G2696,G411);
or gate_637(G2702,G2699,G2701,G374);
and gate_638(G2747,G289,G2728);
and gate_639(G2749,G281,G2728);
and gate_640(G2751,G273,G2728);
and gate_641(G2753,G265,G2728);
and gate_642(G2755,G257,G2728);
and gate_643(G2757,G234,G2741);
and gate_644(G2759,G226,G2741);
and gate_645(G2761,G218,G2741);
and gate_646(G2763,G210,G2741);
and gate_647(G2765,G206,G2741);
not gate_648(G2857,G2847);
or gate_649(G2908,G2906,G2907);
or gate_650(G2911,G2909,G2910);
or gate_651(G2915,G2913,G2914);
or gate_652(G2925,G2922,G2924,G479);
or gate_653(G2930,G2927,G2929,G490);
or gate_654(G2933,G2918,G2920);
or gate_655(G2976,G2973,G2975);
or gate_656(G2985,G2982,G2984);
or gate_657(G2991,G2988,G2990);
or gate_658(G2997,G2994,G2996,G503);
or gate_659(G3004,G3001,G3003,G523);
or gate_660(G3009,G3006,G3008,G534);
or gate_661(G3058,G3056,G3057);
or gate_662(G3062,G3060,G3061);
or gate_663(G3066,G3064,G3065);
or gate_664(G3070,G3068,G3069);
or gate_665(G3076,G3073,G3075,G389);
or gate_666(G3081,G3078,G3080,G400);
or gate_667(G3086,G3083,G3085,G411);
or gate_668(G3091,G3088,G3090,G374);
and gate_669(G3118,G369,G3099);
and gate_670(G3120,G361,G3099);
and gate_671(G3122,G351,G3099);
and gate_672(G3124,G341,G3099);
and gate_673(G3127,G324,G3112);
and gate_674(G3129,G316,G3112);
and gate_675(G3131,G308,G3112);
and gate_676(G3133,G302,G3112);
and gate_677(G3135,G293,G3112);
or gate_678(G3147,G3099,G3126);
and gate_679(G3192,G83,G3187);
and gate_680(G3195,G87,G3187);
and gate_681(G3198,G34,G3187);
and gate_682(G3201,G34,G3187);
or gate_683(G3230,G3228,G3229);
or gate_684(G3236,G3234,G3235);
or gate_685(G3240,G3238,G3239);
or gate_686(G3245,G3243,G3244,G503);
or gate_687(G3251,G3249,G3250,G523);
or gate_688(G3255,G3253,G3254,G534);
or gate_689(G3282,G3280,G3281);
or gate_690(G3285,G3283,G3284);
or gate_691(G3289,G3287,G3288);
or gate_692(G3297,G3295,G3296,G479);
or gate_693(G3301,G3299,G3300,G490);
not gate_694(G3309,G3306);
not gate_695(G3313,G3310);
not gate_696(G3321,G3318);
not gate_697(G3325,G3322);
or gate_698(G3328,G3326,G3327);
and gate_699(G3329,G2405,G446,G3310);
or gate_700(G3335,G3333,G3334);
and gate_701(G3336,G2405,G446,G3322);
and gate_702(G3341,G3555,G3306);
and gate_703(G3345,G3555,G3318);
or gate_704(G3388,G3386,G3387);
or gate_705(G3392,G3390,G3391);
or gate_706(G3396,G3394,G3395);
or gate_707(G3400,G3398,G3399);
or gate_708(G3406,G3403,G3405,G457);
or gate_709(G3411,G3408,G3410,G468);
or gate_710(G3416,G3413,G3415,G422);
or gate_711(G3421,G3418,G3420,G435);
nand gate_712(G3424,G3422,G3423);
nand gate_713(G3433,G3431,G3432);
not gate_714(G3492,G3489);
not gate_715(G3496,G3493);
and gate_716(G3780,G117,G3745,G3757);
and gate_717(G3783,G126,G3745,G3757);
and gate_718(G3786,G127,G3745,G3757);
and gate_719(G3789,G128,G3745,G3757);
and gate_720(G3838,G131,G3803,G3815);
and gate_721(G3841,G129,G3803,G3815);
and gate_722(G3844,G119,G3803,G3815);
and gate_723(G3847,G130,G3803,G3815);
nand gate_724(G3897,G3895,G3896);
nand gate_725(G3906,G3904,G3905);
nand gate_726(G3915,G3913,G3914);
and gate_727(G4011,G122,G3979,G3991);
and gate_728(G4014,G113,G3979,G3991);
and gate_729(G4017,G53,G3979,G3991);
and gate_730(G4020,G114,G3979,G3991);
and gate_731(G4023,G115,G3979,G3991);
and gate_732(G4069,G52,G4037,G4049);
and gate_733(G4072,G112,G4037,G4049);
and gate_734(G4075,G116,G4037,G4049);
and gate_735(G4078,G121,G4037,G4049);
and gate_736(G4081,G123,G4037,G4049);
nand gate_737(G5206,G5116,G5117);
nand gate_738(G5209,G5106,G5107);
and gate_739(G5307,G3233,G3247);
or gate_740(G5322,G3292,G3293);
not gate_741(G5372,G5366);
nand gate_742(G5375,G5366,G5373);
nand gate_743(G5399,G5364,G5365);
not gate_744(G2813,G3015);
or gate_745(G3197,G3195,G3196);
or gate_746(G3200,G3198,G3199);
or gate_747(G3203,G3201,G3202);
or gate_748(G3194,G3192,G3193);
not gate_749(G2570,G2569);
not gate_750(G2576,G2575);
not gate_751(G2582,G2581);
not gate_752(G2588,G2587);
not gate_753(G2664,G2663);
not gate_754(G2670,G2669);
not gate_755(G2676,G2675);
not gate_756(G2682,G2681);
or gate_757(G2767,G2749,G2750);
or gate_758(G2772,G2751,G2752);
or gate_759(G2776,G2753,G2754);
or gate_760(G2780,G2755,G2756);
or gate_761(G2784,G2757,G2758);
or gate_762(G2788,G2759,G2760);
or gate_763(G2794,G2761,G2762);
or gate_764(G2798,G2763,G2764);
or gate_765(G2802,G2765,G2766);
not gate_766(G2912,G2911);
not gate_767(G2916,G2915);
not gate_768(G2936,G2908);
not gate_769(G2977,G2976);
not gate_770(G2986,G2985);
not gate_771(G2992,G2991);
not gate_772(G3059,G3058);
not gate_773(G3063,G3062);
not gate_774(G3067,G3066);
not gate_775(G3071,G3070);
or gate_776(G3137,G3120,G3121);
or gate_777(G3139,G3122,G3123);
or gate_778(G3143,G3124,G3125);
or gate_779(G3151,G3127,G3128);
or gate_780(G3155,G3129,G3130);
or gate_781(G3161,G3131,G3132);
or gate_782(G3165,G3133,G3134);
or gate_783(G3167,G3135,G3136);
not gate_784(G3231,G3230);
not gate_785(G3237,G3236);
not gate_786(G3241,G3240);
not gate_787(G3286,G3285);
not gate_788(G3290,G3289);
and gate_789(G3330,G446,G2382,G3313);
and gate_790(G3337,G446,G2382,G3325);
and gate_791(G3342,G2361,G3309);
and gate_792(G3346,G2361,G3321);
not gate_793(G3348,G3328);
not gate_794(G3352,G3335);
not gate_795(G3389,G3388);
not gate_796(G3393,G3392);
not gate_797(G3397,G3396);
not gate_798(G3401,G3400);
and gate_799(G3845,G3015,G3803,G3823);
or gate_800(G5126,G3118,G3119);
or gate_801(G5178,G2747,G2748);
not gate_802(G5325,G3282);
nand gate_803(G5374,G5369,G5372);
not gate_804(G2810,G2933);
and gate_805(G635,G3197,G3176);
and gate_806(G2878,G24,G2838,G2857);
and gate_807(G2879,G25,G2828,G2857);
and gate_808(G2874,G26,G2838,G2857);
and gate_809(G2875,G81,G2828,G2857);
and gate_810(G703,G3200,G3176);
and gate_811(G2866,G79,G2838,G2857);
and gate_812(G2867,G23,G2828,G2857);
and gate_813(G2870,G82,G2838,G2857);
and gate_814(G2871,G80,G2828,G2857);
and gate_815(G716,G3203,G3176);
and gate_816(G819,G3194,G3176);
and gate_817(G1789,G3147,G514);
and gate_818(G2036,G514,G3147);
and gate_819(G2611,G2570,G2593);
and gate_820(G2615,G2576,G2598);
and gate_821(G2619,G2582,G2603);
and gate_822(G2623,G2588,G2608);
and gate_823(G2705,G2664,G2687);
and gate_824(G2709,G2670,G2692);
and gate_825(G2713,G2676,G2697);
and gate_826(G2717,G2682,G2702);
and gate_827(G2939,G2912,G2925);
and gate_828(G2942,G2916,G2930);
buf gate_829(G2945,G2933);
and gate_830(G3012,G2977,G2997);
and gate_831(G3018,G2986,G3004);
and gate_832(G3021,G2992,G3009);
or gate_833(G3331,G3329,G3330);
or gate_834(G3338,G3336,G3337);
or gate_835(G3343,G3341,G3342,G446);
or gate_836(G3347,G3345,G3346,G446);
not gate_837(G3428,G3424);
not gate_838(G3437,G3433);
and gate_839(G3514,G3433,G3424,G3489);
and gate_840(G3836,G3352,G3803,G3823);
and gate_841(G3852,G3071,G3091);
not gate_842(G5311,G5307);
not gate_843(G3901,G3897);
not gate_844(G3910,G3906);
buf gate_845(G3934,G3915);
buf gate_846(G3938,G3915);
buf gate_847(G4652,G3147);
buf gate_848(G4783,G3147);
buf gate_849(G5137,G3147);
not gate_850(G5212,G5206);
not gate_851(G5213,G5209);
and gate_852(G5260,G3063,G3081);
and gate_853(G5263,G3067,G3086);
and gate_854(G5268,G3401,G3421);
and gate_855(G5271,G3059,G3076);
and gate_856(G5276,G3393,G3411);
and gate_857(G5279,G3397,G3416);
and gate_858(G5289,G3389,G3406);
and gate_859(G5296,G3237,G3251);
and gate_860(G5299,G3241,G3255);
and gate_861(G5304,G3231,G3245);
and gate_862(G5312,G3286,G3297);
and gate_863(G5315,G3290,G3301);
not gate_864(G5328,G5322);
nand gate_865(G5396,G5374,G5375);
not gate_866(G5403,G5399);
and gate_867(G1286,G446,G2802);
not gate_868(G2809,G2936);
not gate_869(G597,G3348);
and gate_870(G1031,G2802,G446);
not gate_871(G636,G635);
or gate_872(G637,G2878,G2879,G2880,G2881);
or gate_873(G671,G2874,G2875,G2876,G2877);
not gate_874(G704,G703);
or gate_875(G705,G2866,G2867,G2868,G2869);
or gate_876(G713,G2870,G2871,G2872,G2873);
not gate_877(G717,G716);
not gate_878(G820,G819);
and gate_879(G1046,G2798,G457);
and gate_880(G1064,G2794,G468);
and gate_881(G1071,G422,G2788);
and gate_882(G1097,G2784,G435);
and gate_883(G1111,G2780,G389);
and gate_884(G1128,G2776,G400);
and gate_885(G1145,G2772,G411);
and gate_886(G1160,G2767,G374);
and gate_887(G1301,G457,G2798);
and gate_888(G1318,G468,G2794);
and gate_889(G1324,G422,G2788);
and gate_890(G1341,G435,G2784);
and gate_891(G1359,G389,G2780);
and gate_892(G1382,G400,G2776);
and gate_893(G1404,G411,G2772);
and gate_894(G1412,G374,G2767);
not gate_895(G1704,G3167);
not gate_896(G1712,G3165);
buf gate_897(G1724,G3165);
and gate_898(G1742,G3161,G479);
and gate_899(G1749,G490,G3155);
and gate_900(G1775,G3151,G503);
and gate_901(G1806,G3143,G523);
and gate_902(G1823,G3139,G534);
not gate_903(G1829,G3137);
buf gate_904(G1837,G3137);
not gate_905(G1958,G3167);
not gate_906(G1966,G3165);
buf gate_907(G1978,G3165);
and gate_908(G1995,G479,G3161);
and gate_909(G2001,G490,G3155);
and gate_910(G2018,G503,G3151);
and gate_911(G2059,G523,G3143);
and gate_912(G2081,G534,G3139);
buf gate_913(G2089,G3137);
not gate_914(G2106,G3137);
buf gate_915(G3170,G3167);
not gate_916(G3332,G3331);
not gate_917(G3339,G3338);
not gate_918(G5132,G5126);
not gate_919(G5184,G5178);
not gate_920(G3853,G3852);
not gate_921(G3874,G3348);
and gate_922(G4076,G2936,G4037,G4056);
buf gate_923(G4116,G2802);
buf gate_924(G4124,G2798);
buf gate_925(G4132,G2794);
buf gate_926(G4140,G2788);
buf gate_927(G4148,G2784);
buf gate_928(G4156,G2780);
buf gate_929(G4164,G2776);
buf gate_930(G4172,G2772);
buf gate_931(G4180,G2767);
nor gate_932(G4228,G422,G2788);
buf gate_933(G4279,G2802);
buf gate_934(G4287,G2798);
buf gate_935(G4295,G2794);
buf gate_936(G4303,G2784);
buf gate_937(G4311,G2780);
buf gate_938(G4319,G2776);
buf gate_939(G4327,G2772);
buf gate_940(G4335,G2788);
buf gate_941(G4343,G2767);
nor gate_942(G4348,G422,G2788);
nor gate_943(G4464,G374,G2767);
buf gate_944(G4628,G3161);
buf gate_945(G4636,G3155);
buf gate_946(G4644,G3151);
buf gate_947(G4660,G3143);
buf gate_948(G4668,G3139);
nor gate_949(G4716,G490,G3155);
buf gate_950(G4767,G3161);
buf gate_951(G4775,G3151);
buf gate_952(G4791,G3143);
buf gate_953(G4799,G3139);
buf gate_954(G4807,G3155);
nor gate_955(G4812,G490,G3155);
buf gate_956(G5118,G3139);
buf gate_957(G5121,G3143);
buf gate_958(G5129,G3137);
buf gate_959(G5134,G3151);
buf gate_960(G5142,G3161);
buf gate_961(G5145,G3155);
buf gate_962(G5152,G3167);
buf gate_963(G5155,G3165);
buf gate_964(G5162,G2788);
buf gate_965(G5165,G2784);
buf gate_966(G5170,G2798);
buf gate_967(G5173,G2794);
buf gate_968(G5181,G2802);
buf gate_969(G5186,G2772);
buf gate_970(G5189,G2767);
buf gate_971(G5196,G2780);
buf gate_972(G5199,G2776);
nand gate_973(G5214,G5209,G5212);
nand gate_974(G5215,G5206,G5213);
not gate_975(G5329,G5325);
nand gate_976(G5330,G5325,G5328);
not gate_977(G2807,G2942);
not gate_978(G2808,G2939);
not gate_979(G2811,G3021);
not gate_980(G2812,G3018);
not gate_981(G2814,G3012);
not gate_982(G2626,G2623);
not gate_983(G2622,G2619);
not gate_984(G2618,G2615);
not gate_985(G2614,G2611);
not gate_986(G2720,G2717);
not gate_987(G2716,G2713);
not gate_988(G2712,G2709);
not gate_989(G2708,G2705);
and gate_990(G639,G637,G2827);
and gate_991(G673,G671,G2827);
and gate_992(G707,G705,G2827);
and gate_993(G715,G713,G2827);
and gate_994(G3731,G2945,G3728,G3721);
not gate_995(G4658,G4652);
nand gate_996(G1777,G4652,G4659);
nand gate_997(G2019,G4783,G4786);
not gate_998(G4787,G4783);
and gate_999(G3350,G3332,G3343);
and gate_1000(G3353,G3339,G3347);
not gate_1001(G5141,G5137);
and gate_1002(G3513,G3428,G3433,G3492);
and gate_1003(G3516,G3424,G3437,G3496);
and gate_1004(G3517,G3437,G3428,G3493);
and gate_1005(G3778,G2717,G3745,G3765);
and gate_1006(G3781,G2713,G3745,G3765);
and gate_1007(G3784,G2709,G3745,G3765);
and gate_1008(G3787,G2705,G3745,G3765);
and gate_1009(G3839,G3021,G3803,G3823);
and gate_1010(G3842,G3018,G3803,G3823);
not gate_1011(G5266,G5260);
not gate_1012(G5267,G5263);
not gate_1013(G5274,G5268);
not gate_1014(G5275,G5271);
not gate_1015(G5302,G5296);
not gate_1016(G5303,G5299);
not gate_1017(G5310,G5304);
nand gate_1018(G3891,G5304,G5311);
not gate_1019(G3937,G3934);
not gate_1020(G3941,G3938);
and gate_1021(G3955,G3906,G3897,G3934);
and gate_1022(G3958,G3910,G3901,G3938);
and gate_1023(G4009,G2623,G3979,G3998);
and gate_1024(G4012,G2619,G3979,G3998);
and gate_1025(G4015,G2615,G3979,G3998);
and gate_1026(G4018,G2611,G3979,G3998);
and gate_1027(G4067,G3012,G4037,G4056);
and gate_1028(G4070,G2942,G4037,G4056);
and gate_1029(G4073,G2939,G4037,G4056);
and gate_1030(G4079,G2945,G4037,G4056);
nand gate_1031(G5239,G5214,G5215);
not gate_1032(G5282,G5276);
not gate_1033(G5283,G5279);
not gate_1034(G5293,G5289);
not gate_1035(G5318,G5312);
not gate_1036(G5319,G5315);
nand gate_1037(G5331,G5322,G5329);
not gate_1038(G5402,G5396);
nand gate_1039(G5405,G5396,G5403);
and gate_1040(G595,G2807,G2808,G2809,G2810);
and gate_1041(G596,G2811,G2812,G2813,G2814);
and gate_1042(G607,G2626,G2622,G2618,G2614);
and gate_1043(G608,G2720,G2716,G2712,G2708);
and gate_1044(G1845,G1704,G1724);
and gate_1045(G1846,G1712,G1704,G1742);
and gate_1046(G2115,G1958,G1978);
and gate_1047(G2116,G1966,G1958,G1995);
not gate_1048(G4122,G4116);
nand gate_1049(G1022,G4116,G4123);
not gate_1050(G4130,G4124);
nand gate_1051(G1033,G4124,G4131);
not gate_1052(G4138,G4132);
nand gate_1053(G1051,G4132,G4139);
not gate_1054(G4146,G4140);
nand gate_1055(G1079,G4140,G4147);
not gate_1056(G4154,G4148);
nand gate_1057(G1088,G4148,G4155);
not gate_1058(G4162,G4156);
nand gate_1059(G1099,G4156,G4163);
not gate_1060(G4170,G4164);
nand gate_1061(G1115,G4164,G4171);
not gate_1062(G4178,G4172);
nand gate_1063(G1133,G4172,G4179);
not gate_1064(G4186,G4180);
nand gate_1065(G1151,G4180,G4187);
not gate_1066(G4234,G4228);
nand gate_1067(G1276,G4279,G4282);
not gate_1068(G4283,G4279);
nand gate_1069(G1287,G4287,G4290);
not gate_1070(G4291,G4287);
nand gate_1071(G1305,G4295,G4298);
not gate_1072(G4299,G4295);
nand gate_1073(G1330,G4303,G4306);
not gate_1074(G4307,G4303);
nand gate_1075(G1342,G4311,G4314);
not gate_1076(G4315,G4311);
nand gate_1077(G1363,G4319,G4322);
not gate_1078(G4323,G4319);
nand gate_1079(G1388,G4327,G4330);
not gate_1080(G4331,G4327);
nand gate_1081(G1420,G4335,G4338);
not gate_1082(G4339,G4335);
nand gate_1083(G1428,G4343,G4346);
not gate_1084(G4347,G4343);
not gate_1085(G4634,G4628);
nand gate_1086(G1729,G4628,G4635);
not gate_1087(G4642,G4636);
nand gate_1088(G1757,G4636,G4643);
not gate_1089(G4650,G4644);
nand gate_1090(G1766,G4644,G4651);
nand gate_1091(G1776,G4655,G4658);
not gate_1092(G4666,G4660);
nand gate_1093(G1793,G4660,G4667);
not gate_1094(G4674,G4668);
nand gate_1095(G1811,G4668,G4675);
and gate_1096(G1849,G1712,G1742);
and gate_1097(G1852,G1712,G1742);
and gate_1098(G1875,G54,G1829);
not gate_1099(G4722,G4716);
nand gate_1100(G1982,G4767,G4770);
not gate_1101(G4771,G4767);
nand gate_1102(G2007,G4775,G4778);
not gate_1103(G4779,G4775);
nand gate_1104(G2020,G4780,G4787);
nand gate_1105(G2040,G4791,G4794);
not gate_1106(G4795,G4791);
nand gate_1107(G2065,G4799,G4802);
not gate_1108(G4803,G4799);
nand gate_1109(G2097,G4807,G4810);
not gate_1110(G4811,G4807);
and gate_1111(G2119,G1966,G1995);
and gate_1112(G2122,G1966,G1995);
not gate_1113(G5124,G5118);
not gate_1114(G5125,G5121);
nand gate_1115(G3452,G5129,G5132);
not gate_1116(G5133,G5129);
not gate_1117(G5140,G5134);
nand gate_1118(G3462,G5134,G5141);
not gate_1119(G5168,G5162);
not gate_1120(G5169,G5165);
not gate_1121(G5176,G5170);
not gate_1122(G5177,G5173);
nand gate_1123(G3484,G5181,G5184);
not gate_1124(G5185,G5181);
nor gate_1125(G3515,G3513,G3514);
nor gate_1126(G3518,G3516,G3517);
not gate_1127(G3857,G3853);
nand gate_1128(G3860,G5263,G5266);
nand gate_1129(G3861,G5260,G5267);
nand gate_1130(G3869,G5271,G5274);
nand gate_1131(G3870,G5268,G5275);
not gate_1132(G3878,G3874);
nand gate_1133(G3881,G5299,G5302);
nand gate_1134(G3882,G5296,G5303);
nand gate_1135(G3890,G5307,G5310);
and gate_1136(G3954,G3901,G3906,G3937);
and gate_1137(G3957,G3897,G3910,G3941);
and gate_1138(G4021,G3353,G3979,G3998);
not gate_1139(G4099,G3170);
buf gate_1140(G4236,G1071);
not gate_1141(G4354,G4348);
buf gate_1142(G4406,G1324);
not gate_1143(G4470,G4464);
buf gate_1144(G4552,G1412);
buf gate_1145(G4679,G1829);
buf gate_1146(G4687,G1704);
buf gate_1147(G4695,G1704);
buf gate_1148(G4703,G1712);
buf gate_1149(G4711,G1712);
buf gate_1150(G4724,G1749);
not gate_1151(G4818,G4812);
buf gate_1152(G4855,G1958);
buf gate_1153(G4865,G1966);
buf gate_1154(G4870,G2001);
buf gate_1155(G4913,G1958);
buf gate_1156(G4923,G1966);
buf gate_1157(G4951,G2106);
buf gate_1158(G5006,G2089);
buf gate_1159(G5039,G2106);
not gate_1160(G5148,G5142);
not gate_1161(G5149,G5145);
not gate_1162(G5158,G5152);
not gate_1163(G5159,G5155);
not gate_1164(G5192,G5186);
not gate_1165(G5193,G5189);
not gate_1166(G5202,G5196);
not gate_1167(G5203,G5199);
nand gate_1168(G5284,G5279,G5282);
nand gate_1169(G5285,G5276,G5283);
nand gate_1170(G5320,G5315,G5318);
nand gate_1171(G5321,G5312,G5319);
nand gate_1172(G5386,G5330,G5331);
nand gate_1173(G5404,G5399,G5402);
and gate_1174(G598,G595,G596,G597);
not gate_1175(G609,G3350);
nand gate_1176(G1021,G4119,G4122);
nand gate_1177(G1032,G4127,G4130);
nand gate_1178(G1050,G4135,G4138);
nand gate_1179(G1078,G4143,G4146);
nand gate_1180(G1087,G4151,G4154);
nand gate_1181(G1098,G4159,G4162);
nand gate_1182(G1114,G4167,G4170);
nand gate_1183(G1132,G4175,G4178);
nand gate_1184(G1150,G4183,G4186);
nand gate_1185(G1277,G4276,G4283);
nand gate_1186(G1288,G4284,G4291);
nand gate_1187(G1306,G4292,G4299);
nand gate_1188(G1331,G4300,G4307);
nand gate_1189(G1343,G4308,G4315);
nand gate_1190(G1364,G4316,G4323);
nand gate_1191(G1389,G4324,G4331);
nand gate_1192(G1421,G4332,G4339);
nand gate_1193(G1429,G4340,G4347);
nand gate_1194(G1728,G4631,G4634);
nand gate_1195(G1756,G4639,G4642);
nand gate_1196(G1765,G4647,G4650);
nand gate_1197(G1778,G1776,G1777);
nand gate_1198(G1792,G4663,G4666);
nand gate_1199(G1810,G4671,G4674);
nand gate_1200(G1983,G4764,G4771);
nand gate_1201(G2008,G4772,G4779);
nand gate_1202(G2021,G2019,G2020);
nand gate_1203(G2041,G4788,G4795);
nand gate_1204(G2066,G4796,G4803);
nand gate_1205(G2098,G4804,G4811);
nand gate_1206(G3443,G5121,G5124);
nand gate_1207(G3444,G5118,G5125);
nand gate_1208(G3453,G5126,G5133);
nand gate_1209(G3461,G5137,G5140);
nand gate_1210(G3466,G5165,G5168);
nand gate_1211(G3467,G5162,G5169);
nand gate_1212(G3475,G5173,G5176);
nand gate_1213(G3476,G5170,G5177);
nand gate_1214(G3485,G5178,G5185);
not gate_1215(G5243,G5239);
nand gate_1216(G3862,G3860,G3861);
nand gate_1217(G3871,G3869,G3870);
nand gate_1218(G3883,G3881,G3882);
nand gate_1219(G3892,G3890,G3891);
nor gate_1220(G3956,G3954,G3955);
nor gate_1221(G3959,G3957,G3958);
or gate_1222(G4756,G1837,G1875);
nand gate_1223(G5150,G5145,G5148);
nand gate_1224(G5151,G5142,G5149);
nand gate_1225(G5160,G5155,G5158);
nand gate_1226(G5161,G5152,G5159);
nand gate_1227(G5194,G5189,G5192);
nand gate_1228(G5195,G5186,G5193);
nand gate_1229(G5204,G5199,G5202);
nand gate_1230(G5205,G5196,G5203);
nand gate_1231(G5236,G3518,G3515);
buf gate_1232(G5286,G3350);
nand gate_1233(G5379,G5284,G5285);
nand gate_1234(G5389,G5320,G5321);
nand gate_1235(G5425,G5404,G5405);
and gate_1236(G610,G607,G608,G609);
nand gate_1237(G1023,G1021,G1022);
nand gate_1238(G1034,G1032,G1033);
nand gate_1239(G1052,G1050,G1051);
nand gate_1240(G1080,G1078,G1079);
nand gate_1241(G1089,G1087,G1088);
nand gate_1242(G1100,G1098,G1099);
nand gate_1243(G1116,G1114,G1115);
nand gate_1244(G1134,G1132,G1133);
nand gate_1245(G1152,G1150,G1151);
not gate_1246(G4242,G4236);
nand gate_1247(G1278,G1276,G1277);
nand gate_1248(G1289,G1287,G1288);
nand gate_1249(G1307,G1305,G1306);
nand gate_1250(G1332,G1330,G1331);
nand gate_1251(G1344,G1342,G1343);
nand gate_1252(G1365,G1363,G1364);
nand gate_1253(G1390,G1388,G1389);
nand gate_1254(G1422,G1420,G1421);
nand gate_1255(G1430,G1428,G1429);
nand gate_1256(G1730,G1728,G1729);
nand gate_1257(G1758,G1756,G1757);
nand gate_1258(G1767,G1765,G1766);
nand gate_1259(G1794,G1792,G1793);
nand gate_1260(G1812,G1810,G1811);
nand gate_1261(G1876,G4679,G4682);
not gate_1262(G4683,G4679);
not gate_1263(G4691,G4687);
not gate_1264(G4699,G4695);
not gate_1265(G4707,G4703);
not gate_1266(G4715,G4711);
not gate_1267(G4730,G4724);
nand gate_1268(G1984,G1982,G1983);
nand gate_1269(G2009,G2007,G2008);
nand gate_1270(G2042,G2040,G2041);
nand gate_1271(G2067,G2065,G2066);
nand gate_1272(G2099,G2097,G2098);
not gate_1273(G4869,G4865);
not gate_1274(G4927,G4923);
nand gate_1275(G3445,G3443,G3444);
nand gate_1276(G3454,G3452,G3453);
nand gate_1277(G3463,G3461,G3462);
nand gate_1278(G3468,G3466,G3467);
nand gate_1279(G3477,G3475,G3476);
nand gate_1280(G3486,G3484,G3485);
and gate_1281(G4103,G4099,G3170);
not gate_1282(G4412,G4406);
not gate_1283(G4558,G4552);
not gate_1284(G4859,G4855);
not gate_1285(G4876,G4870);
not gate_1286(G4917,G4913);
not gate_1287(G4955,G4951);
not gate_1288(G5012,G5006);
not gate_1289(G5043,G5039);
nand gate_1290(G5216,G5160,G5161);
nand gate_1291(G5219,G5150,G5151);
nand gate_1292(G5226,G5204,G5205);
nand gate_1293(G5229,G5194,G5195);
not gate_1294(G5392,G5386);
nand gate_1295(G5422,G3959,G3956);
and gate_1296(G1866,G1778,G1806);
nand gate_1297(G1877,G4676,G4683);
not gate_1298(G4762,G4756);
and gate_1299(G2142,G2021,G2059);
and gate_1300(G2146,G2021,G2059);
not gate_1301(G5242,G5236);
nand gate_1302(G3532,G5236,G5243);
not gate_1303(G3866,G3862);
not gate_1304(G3887,G3883);
buf gate_1305(G3918,G3871);
buf gate_1306(G3922,G3871);
buf gate_1307(G3926,G3892);
buf gate_1308(G3930,G3892);
not gate_1309(G5429,G5425);
or gate_1310(G4104,G4099,G4103);
buf gate_1311(G4743,G1778);
buf gate_1312(G4991,G2021);
buf gate_1313(G5001,G2021);
not gate_1314(G5292,G5286);
nand gate_1315(G5295,G5286,G5293);
not gate_1316(G5383,G5379);
not gate_1317(G5393,G5389);
nand gate_1318(G5394,G5389,G5392);
and gate_1319(G1439,G1278,G1301);
and gate_1320(G1440,G1289,G1278,G1318);
and gate_1321(G1441,G1307,G1278,G1324,G1289);
and gate_1322(G1847,G1730,G1704,G1749,G1712);
and gate_1323(G1168,G1023,G1046);
and gate_1324(G1169,G1034,G1023,G1064);
and gate_1325(G1170,G1052,G1023,G1071,G1034);
and gate_1326(G2117,G1984,G1958,G2001,G1966);
not gate_1327(G1086,G1080);
and gate_1328(G1166,G1034,G1080,G1052,G1023);
and gate_1329(G1171,G1034,G1064);
and gate_1330(G1172,G1052,G1071,G1034);
and gate_1331(G1173,G1080,G1052,G1034);
and gate_1332(G1174,G1034,G1064);
and gate_1333(G1175,G1071,G1052,G1034);
and gate_1334(G1176,G1052,G1071);
and gate_1335(G1177,G1080,G1052);
and gate_1336(G1178,G1052,G1071);
and gate_1337(G1179,G1100,G1152,G1116,G1089,G1134);
and gate_1338(G1181,G1089,G1111);
and gate_1339(G1182,G1100,G1089,G1128);
and gate_1340(G1183,G1116,G1089,G1145,G1100);
and gate_1341(G1184,G1134,G1116,G1089,G1160,G1100);
and gate_1342(G1188,G1100,G1128);
and gate_1343(G1189,G1116,G1145,G1100);
and gate_1344(G1190,G1134,G1116,G1160,G1100);
and gate_1345(G1191,G4,G1152,G1116,G1134,G1100);
and gate_1346(G1192,G1145,G1116);
and gate_1347(G1193,G1134,G1116,G1160);
and gate_1348(G1194,G4,G1152,G1116,G1134);
and gate_1349(G1195,G1134,G1160);
and gate_1350(G1196,G4,G1152,G1134);
and gate_1351(G1197,G4,G1152);
and gate_1352(G1437,G1422,G1307,G1289,G1278);
and gate_1353(G1442,G1289,G1318);
and gate_1354(G1443,G1307,G1324,G1289);
and gate_1355(G1444,G1422,G1307,G1289);
and gate_1356(G1445,G1289,G1318);
and gate_1357(G1446,G1307,G1324,G1289);
and gate_1358(G1447,G1307,G1324);
and gate_1359(G1451,G1430,G1390,G1365,G1344,G1332);
and gate_1360(G1454,G1332,G1359);
and gate_1361(G1455,G1344,G1332,G1382);
and gate_1362(G1456,G1365,G1332,G1404,G1344);
and gate_1363(G1457,G1390,G1365,G1332,G1412,G1344);
and gate_1364(G1465,G1344,G1382);
and gate_1365(G1466,G1365,G1404,G1344);
and gate_1366(G1467,G1390,G1365,G1412,G1344);
and gate_1367(G1468,G1430,G1365,G1344,G1390);
and gate_1368(G1469,G1344,G1382);
and gate_1369(G1470,G1365,G1404,G1344);
and gate_1370(G1471,G1390,G1365,G1412,G1344);
and gate_1371(G1472,G1365,G1404);
and gate_1372(G1473,G1390,G1365,G1412);
and gate_1373(G1474,G1430,G1365,G1390);
and gate_1374(G1475,G1365,G1404);
and gate_1375(G1476,G1390,G1365,G1412);
and gate_1376(G1477,G1390,G1412);
and gate_1377(G1481,G1422,G1307);
and gate_1378(G1482,G1430,G1390);
not gate_1379(G1764,G1758);
and gate_1380(G1843,G1712,G1758,G1730,G1704);
and gate_1381(G1850,G1730,G1749,G1712);
and gate_1382(G1851,G1758,G1730,G1712);
and gate_1383(G1853,G1749,G1730,G1712);
and gate_1384(G1854,G1730,G1749);
and gate_1385(G1855,G1758,G1730);
and gate_1386(G1856,G1730,G1749);
and gate_1387(G1857,G1778,G1829,G1794,G1767,G1812);
and gate_1388(G1859,G1767,G1789);
and gate_1389(G1860,G1778,G1767,G1806);
and gate_1390(G1861,G1794,G1767,G1823,G1778);
and gate_1391(G1862,G1812,G1794,G1767,G1837,G1778);
and gate_1392(G1867,G1794,G1823,G1778);
and gate_1393(G1868,G1812,G1794,G1837,G1778);
and gate_1394(G1869,G54,G1829,G1794,G1812,G1778);
and gate_1395(G1870,G1823,G1794);
and gate_1396(G1871,G1812,G1794,G1837);
and gate_1397(G1872,G54,G1829,G1794,G1812);
and gate_1398(G1873,G1812,G1837);
and gate_1399(G1874,G54,G1829,G1812);
nand gate_1400(G1878,G1876,G1877);
and gate_1401(G2113,G2099,G1984,G1966,G1958);
and gate_1402(G2120,G1984,G2001,G1966);
and gate_1403(G2121,G2099,G1984,G1966);
and gate_1404(G2123,G1984,G2001,G1966);
and gate_1405(G2124,G1984,G2001);
and gate_1406(G2128,G2106,G2067,G2042,G2021,G2009);
and gate_1407(G2131,G2009,G2036);
and gate_1408(G2132,G2021,G2009,G2059);
and gate_1409(G2133,G2042,G2009,G2081,G2021);
and gate_1410(G2134,G2067,G2042,G2009,G2089,G2021);
and gate_1411(G2143,G2042,G2081,G2021);
and gate_1412(G2144,G2067,G2042,G2089,G2021);
and gate_1413(G2145,G2106,G2042,G2021,G2067);
and gate_1414(G2147,G2042,G2081,G2021);
and gate_1415(G2148,G2067,G2042,G2089,G2021);
and gate_1416(G2149,G2042,G2081);
and gate_1417(G2150,G2067,G2042,G2089);
and gate_1418(G2151,G2106,G2042,G2067);
and gate_1419(G2152,G2042,G2081);
and gate_1420(G2153,G2067,G2042,G2089);
and gate_1421(G2154,G2067,G2089);
and gate_1422(G2158,G2099,G1984);
and gate_1423(G2159,G2106,G2067);
not gate_1424(G3449,G3445);
not gate_1425(G3458,G3454);
not gate_1426(G3472,G3468);
not gate_1427(G3481,G3477);
buf gate_1428(G3497,G3463);
buf gate_1429(G3501,G3463);
buf gate_1430(G3505,G3486);
buf gate_1431(G3509,G3486);
nand gate_1432(G3531,G5239,G5242);
not gate_1433(G5428,G5422);
nand gate_1434(G3967,G5422,G5429);
buf gate_1435(G4191,G1152);
buf gate_1436(G4199,G1023);
buf gate_1437(G4207,G1023);
buf gate_1438(G4215,G1034);
buf gate_1439(G4223,G1034);
buf gate_1440(G4231,G1052);
buf gate_1441(G4239,G1052);
buf gate_1442(G4247,G1089);
buf gate_1443(G4255,G1100);
buf gate_1444(G4263,G1116);
buf gate_1445(G4271,G1134);
buf gate_1446(G4371,G1422);
buf gate_1447(G4381,G1307);
buf gate_1448(G4391,G1278);
buf gate_1449(G4401,G1289);
buf gate_1450(G4429,G1422);
buf gate_1451(G4439,G1307);
buf gate_1452(G4449,G1278);
buf gate_1453(G4459,G1289);
buf gate_1454(G4497,G1430);
buf gate_1455(G4507,G1390);
buf gate_1456(G4517,G1332);
buf gate_1457(G4527,G1365);
buf gate_1458(G4537,G1344);
buf gate_1459(G4547,G1344);
buf gate_1460(G4585,G1430);
buf gate_1461(G4595,G1390);
buf gate_1462(G4605,G1332);
buf gate_1463(G4615,G1365);
buf gate_1464(G4719,G1730);
buf gate_1465(G4727,G1730);
buf gate_1466(G4735,G1767);
buf gate_1467(G4751,G1794);
buf gate_1468(G4759,G1812);
buf gate_1469(G4835,G2099);
buf gate_1470(G4845,G1984);
buf gate_1471(G4893,G2099);
buf gate_1472(G4903,G1984);
buf gate_1473(G4961,G2067);
buf gate_1474(G4971,G2009);
buf gate_1475(G4981,G2042);
buf gate_1476(G5049,G2067);
buf gate_1477(G5059,G2009);
buf gate_1478(G5069,G2042);
not gate_1479(G5222,G5216);
not gate_1480(G5223,G5219);
not gate_1481(G5232,G5226);
not gate_1482(G5233,G5229);
nand gate_1483(G5294,G5289,G5292);
nand gate_1484(G5395,G5386,G5393);
or gate_1485(G589,G1286,G1439,G1440,G1441);
or gate_1486(G616,G3167,G1845,G1846,G1847);
or gate_1487(G619,G1031,G1168,G1169,G1170);
or gate_1488(G627,G3167,G2115,G2116,G2117);
or gate_1489(G1185,G1097,G1181,G1182,G1183,G1184);
or gate_1490(G1448,G1318,G1447);
or gate_1491(G1458,G1341,G1454,G1455,G1456,G1457);
or gate_1492(G1478,G1404,G1477);
or gate_1493(G1863,G1775,G1859,G1860,G1861,G1862);
not gate_1494(G4747,G4743);
or gate_1495(G2125,G1995,G2124);
or gate_1496(G2135,G2018,G2131,G2132,G2133,G2134);
or gate_1497(G2155,G2081,G2154);
not gate_1498(G4995,G4991);
not gate_1499(G5005,G5001);
nand gate_1500(G3533,G3531,G3532);
not gate_1501(G3921,G3918);
not gate_1502(G3925,G3922);
not gate_1503(G3929,G3926);
not gate_1504(G3933,G3930);
and gate_1505(G3943,G3862,G3853,G3918);
and gate_1506(G3946,G3866,G3857,G3922);
and gate_1507(G3949,G3883,G3874,G3926);
and gate_1508(G3952,G3887,G3878,G3930);
nand gate_1509(G3966,G5425,G5428);
nand gate_1510(G4107,G4104,G132);
or gate_1511(G4196,G1046,G1171,G1172,G1173);
nor gate_1512(G4204,G1046,G1174,G1175);
or gate_1513(G4212,G1064,G1176,G1177);
nor gate_1514(G4220,G1064,G1178);
or gate_1515(G4244,G1111,G1188,G1189,G1190,G1191);
or gate_1516(G4252,G1128,G1192,G1193,G1194);
or gate_1517(G4260,G1145,G1195,G1196);
or gate_1518(G4268,G1160,G1197);
or gate_1519(G4361,G1301,G1442,G1443,G1444);
nor gate_1520(G4419,G1301,G1445,G1446);
or gate_1521(G4467,G1382,G1472,G1473,G1474);
or gate_1522(G4487,G1359,G1465,G1466,G1467,G1468);
nor gate_1523(G4555,G1382,G1475,G1476);
nor gate_1524(G4575,G1359,G1469,G1470,G1471);
or gate_1525(G4684,G1724,G1849,G1850,G1851);
nor gate_1526(G4692,G1724,G1852,G1853);
or gate_1527(G4700,G1742,G1854,G1855);
nor gate_1528(G4708,G1742,G1856);
or gate_1529(G4732,G1789,G1866,G1867,G1868,G1869);
or gate_1530(G4740,G1806,G1870,G1871,G1872);
or gate_1531(G4748,G1823,G1873,G1874);
or gate_1532(G4825,G1978,G2119,G2120,G2121);
nor gate_1533(G4883,G1978,G2122,G2123);
or gate_1534(G4928,G2059,G2149,G2150,G2151);
or gate_1535(G4941,G2036,G2142,G2143,G2144,G2145);
nor gate_1536(G5009,G2059,G2152,G2153);
nor gate_1537(G5029,G2036,G2146,G2147,G2148);
nand gate_1538(G5224,G5219,G5222);
nand gate_1539(G5225,G5216,G5223);
nand gate_1540(G5234,G5229,G5232);
nand gate_1541(G5235,G5226,G5233);
nand gate_1542(G5376,G5294,G5295);
nand gate_1543(G5417,G5394,G5395);
not gate_1544(G576,G1878);
and gate_1545(G588,G1437,G1451);
and gate_1546(G615,G1843,G1857);
and gate_1547(G626,G2113,G2128);
and gate_1548(G632,G1166,G1179);
nand gate_1549(G1198,G4191,G4194);
not gate_1550(G4195,G4191);
not gate_1551(G4203,G4199);
not gate_1552(G4211,G4207);
not gate_1553(G4219,G4215);
not gate_1554(G4227,G4223);
nand gate_1555(G1217,G4231,G4234);
not gate_1556(G4235,G4231);
nand gate_1557(G1221,G4239,G4242);
not gate_1558(G4243,G4239);
and gate_1559(G1224,G1179,G4);
not gate_1560(G4251,G4247);
not gate_1561(G4259,G4255);
not gate_1562(G4267,G4263);
not gate_1563(G4275,G4271);
not gate_1564(G1453,G1451);
not gate_1565(G4405,G4401);
not gate_1566(G4463,G4459);
not gate_1567(G4541,G4537);
not gate_1568(G4551,G4547);
nand gate_1569(G1895,G4719,G4722);
not gate_1570(G4723,G4719);
nand gate_1571(G1899,G4727,G4730);
not gate_1572(G4731,G4727);
and gate_1573(G1902,G1857,G54);
not gate_1574(G4739,G4735);
not gate_1575(G4755,G4751);
nand gate_1576(G1929,G4759,G4762);
not gate_1577(G4763,G4759);
not gate_1578(G2130,G2128);
not gate_1579(G3500,G3497);
not gate_1580(G3504,G3501);
not gate_1581(G3508,G3505);
not gate_1582(G3512,G3509);
and gate_1583(G3520,G3454,G3445,G3497);
and gate_1584(G3523,G3458,G3449,G3501);
and gate_1585(G3526,G3477,G3468,G3505);
and gate_1586(G3529,G3481,G3472,G3509);
buf gate_1587(G1002,G3533);
and gate_1588(G3837,G1878,G3795,G3823);
and gate_1589(G3942,G3857,G3862,G3921);
and gate_1590(G3945,G3853,G3866,G3925);
and gate_1591(G3948,G3878,G3883,G3929);
and gate_1592(G3951,G3874,G3887,G3933);
nand gate_1593(G3968,G3966,G3967);
not gate_1594(G4375,G4371);
not gate_1595(G4385,G4381);
not gate_1596(G4395,G4391);
not gate_1597(G4433,G4429);
not gate_1598(G4443,G4439);
not gate_1599(G4453,G4449);
not gate_1600(G4501,G4497);
not gate_1601(G4511,G4507);
not gate_1602(G4521,G4517);
not gate_1603(G4531,G4527);
not gate_1604(G4619,G4615);
not gate_1605(G4589,G4585);
not gate_1606(G4599,G4595);
not gate_1607(G4609,G4605);
not gate_1608(G4839,G4835);
not gate_1609(G4849,G4845);
not gate_1610(G4897,G4893);
not gate_1611(G4907,G4903);
not gate_1612(G4965,G4961);
not gate_1613(G4975,G4971);
not gate_1614(G4985,G4981);
not gate_1615(G5073,G5069);
not gate_1616(G5053,G5049);
not gate_1617(G5063,G5059);
nand gate_1618(G5247,G5224,G5225);
nand gate_1619(G5255,G5234,G5235);
and gate_1620(G590,G1437,G1458);
and gate_1621(G617,G1863,G1843);
and gate_1622(G620,G1185,G1166);
and gate_1623(G628,G2113,G2135);
not gate_1624(G3535,G3533);
nand gate_1625(G1199,G4188,G4195);
not gate_1626(G4202,G4196);
nand gate_1627(G1204,G4196,G4203);
not gate_1628(G4210,G4204);
nand gate_1629(G1207,G4204,G4211);
not gate_1630(G4218,G4212);
nand gate_1631(G1211,G4212,G4219);
not gate_1632(G4226,G4220);
nand gate_1633(G1214,G4220,G4227);
nand gate_1634(G1218,G4228,G4235);
nand gate_1635(G1222,G4236,G4243);
or gate_1636(G1225,G1185,G1224);
not gate_1637(G4250,G4244);
nand gate_1638(G1237,G4244,G4251);
not gate_1639(G4258,G4252);
nand gate_1640(G1242,G4252,G4259);
not gate_1641(G4266,G4260);
nand gate_1642(G1247,G4260,G4267);
not gate_1643(G4274,G4268);
nand gate_1644(G1252,G4268,G4275);
not gate_1645(G1462,G1458);
not gate_1646(G4690,G4684);
nand gate_1647(G1882,G4684,G4691);
not gate_1648(G4698,G4692);
nand gate_1649(G1885,G4692,G4699);
not gate_1650(G4706,G4700);
nand gate_1651(G1889,G4700,G4707);
not gate_1652(G4714,G4708);
nand gate_1653(G1892,G4708,G4715);
nand gate_1654(G1896,G4716,G4723);
nand gate_1655(G1900,G4724,G4731);
or gate_1656(G1903,G1863,G1902);
not gate_1657(G4738,G4732);
nand gate_1658(G1915,G4732,G4739);
not gate_1659(G4746,G4740);
nand gate_1660(G1920,G4740,G4747);
not gate_1661(G4754,G4748);
nand gate_1662(G1925,G4748,G4755);
nand gate_1663(G1930,G4756,G4763);
not gate_1664(G2139,G2135);
and gate_1665(G3519,G3449,G3454,G3500);
and gate_1666(G3522,G3445,G3458,G3504);
and gate_1667(G3525,G3472,G3477,G3508);
and gate_1668(G3528,G3468,G3481,G3512);
or gate_1669(G3848,G3836,G3837,G3838);
nor gate_1670(G3944,G3942,G3943);
nor gate_1671(G3947,G3945,G3946);
nor gate_1672(G3950,G3948,G3949);
nor gate_1673(G3953,G3951,G3952);
not gate_1674(G5421,G5417);
buf gate_1675(G1004,G3968);
and gate_1676(G4111,G4104,G4107);
and gate_1677(G4112,G4107,G132);
or gate_1678(G4351,G1448,G1481);
not gate_1679(G4365,G4361);
not gate_1680(G4409,G1448);
not gate_1681(G4423,G4419);
not gate_1682(G4471,G4467);
nand gate_1683(G4472,G4467,G4470);
or gate_1684(G4477,G1478,G1482);
not gate_1685(G4491,G4487);
not gate_1686(G4559,G4555);
nand gate_1687(G4560,G4555,G4558);
not gate_1688(G4565,G1478);
not gate_1689(G4579,G4575);
or gate_1690(G4815,G2125,G2158);
not gate_1691(G4829,G4825);
not gate_1692(G4873,G2125);
not gate_1693(G4887,G4883);
or gate_1694(G4931,G2155,G2159);
not gate_1695(G4934,G4928);
not gate_1696(G4945,G4941);
not gate_1697(G5013,G5009);
nand gate_1698(G5014,G5009,G5012);
not gate_1699(G5019,G2155);
not gate_1700(G5033,G5029);
not gate_1701(G5382,G5376);
nand gate_1702(G5385,G5376,G5383);
or gate_1703(G591,G589,G590);
or gate_1704(G618,G616,G617);
or gate_1705(G621,G619,G620);
or gate_1706(G629,G627,G628);
not gate_1707(G3970,G3968);
nand gate_1708(G1200,G1198,G1199);
nand gate_1709(G1203,G4199,G4202);
nand gate_1710(G1206,G4207,G4210);
nand gate_1711(G1210,G4215,G4218);
nand gate_1712(G1213,G4223,G4226);
nand gate_1713(G1219,G1217,G1218);
nand gate_1714(G1223,G1221,G1222);
nand gate_1715(G1236,G4247,G4250);
nand gate_1716(G1241,G4255,G4258);
nand gate_1717(G1246,G4263,G4266);
nand gate_1718(G1251,G4271,G4274);
nand gate_1719(G1881,G4687,G4690);
nand gate_1720(G1884,G4695,G4698);
nand gate_1721(G1888,G4703,G4706);
nand gate_1722(G1891,G4711,G4714);
nand gate_1723(G1897,G1895,G1896);
nand gate_1724(G1901,G1899,G1900);
nand gate_1725(G1914,G4735,G4738);
nand gate_1726(G1919,G4743,G4746);
nand gate_1727(G1924,G4751,G4754);
nand gate_1728(G1931,G1929,G1930);
nor gate_1729(G3521,G3519,G3520);
nor gate_1730(G3524,G3522,G3523);
nor gate_1731(G3527,G3525,G3526);
nor gate_1732(G3530,G3528,G3529);
not gate_1733(G5251,G5247);
not gate_1734(G5259,G5255);
or gate_1735(G4113,G4111,G4112);
nand gate_1736(G4473,G4464,G4471);
nand gate_1737(G4561,G4552,G4559);
nand gate_1738(G5015,G5006,G5013);
nand gate_1739(G5384,G5379,G5382);
nand gate_1740(G5406,G3947,G3944);
nand gate_1741(G5414,G3953,G3950);
and gate_1742(G1664,G3848,G1621,G1645);
and gate_1743(G2335,G3848,G2293,G2316);
and gate_1744(G718,G3848,G2430,G2454);
not gate_1745(G822,G3848);
and gate_1746(G855,G3848,G2488,G2512);
nand gate_1747(G1205,G1203,G1204);
nand gate_1748(G1208,G1206,G1207);
nand gate_1749(G1212,G1210,G1211);
nand gate_1750(G1215,G1213,G1214);
not gate_1751(G1220,G1219);
not gate_1752(G1231,G1225);
nand gate_1753(G1238,G1236,G1237);
nand gate_1754(G1243,G1241,G1242);
nand gate_1755(G1248,G1246,G1247);
nand gate_1756(G1253,G1251,G1252);
and gate_1757(G1272,G1225,G1086);
and gate_1758(G1483,G1462,G1453);
nand gate_1759(G1883,G1881,G1882);
nand gate_1760(G1886,G1884,G1885);
nand gate_1761(G1890,G1888,G1889);
nand gate_1762(G1893,G1891,G1892);
not gate_1763(G1898,G1897);
not gate_1764(G1909,G1903);
nand gate_1765(G1916,G1914,G1915);
nand gate_1766(G1921,G1919,G1920);
nand gate_1767(G1926,G1924,G1925);
and gate_1768(G1953,G1903,G1764);
and gate_1769(G2160,G2139,G2130);
not gate_1770(G4355,G4351);
nand gate_1771(G4356,G4351,G4354);
not gate_1772(G4413,G4409);
nand gate_1773(G4414,G4409,G4412);
nand gate_1774(G4474,G4472,G4473);
not gate_1775(G4481,G4477);
nand gate_1776(G4562,G4560,G4561);
not gate_1777(G4569,G4565);
not gate_1778(G4819,G4815);
nand gate_1779(G4820,G4815,G4818);
not gate_1780(G4877,G4873);
nand gate_1781(G4878,G4873,G4876);
not gate_1782(G4935,G4931);
nand gate_1783(G4936,G4931,G4934);
nand gate_1784(G5016,G5014,G5015);
not gate_1785(G5023,G5019);
nand gate_1786(G5244,G3524,G3521);
nand gate_1787(G5252,G3530,G3527);
nand gate_1788(G5409,G5384,G5385);
not gate_1789(G566,G1200);
not gate_1790(G577,G1931);
and gate_1791(G3733,G4113,G3724,G3721);
not gate_1792(G1209,G1208);
not gate_1793(G1216,G1215);
and gate_1794(G1257,G1225,G1205);
and gate_1795(G1262,G1225,G1212);
and gate_1796(G1267,G1225,G1220);
not gate_1797(G1887,G1886);
not gate_1798(G1894,G1893);
and gate_1799(G1935,G1903,G1883);
and gate_1800(G1943,G1903,G1890);
and gate_1801(G1948,G1903,G1898);
and gate_1802(G3779,G1200,G3737,G3765);
and gate_1803(G3840,G1931,G3795,G3823);
not gate_1804(G5412,G5406);
not gate_1805(G5420,G5414);
nand gate_1806(G3964,G5414,G5421);
nand gate_1807(G4357,G4348,G4355);
nand gate_1808(G4415,G4406,G4413);
nand gate_1809(G4821,G4812,G4819);
nand gate_1810(G4879,G4870,G4877);
nand gate_1811(G4937,G4928,G4935);
not gate_1812(G567,G1253);
not gate_1813(G568,G1248);
not gate_1814(G569,G1243);
not gate_1815(G570,G1238);
not gate_1816(G578,G1926);
not gate_1817(G579,G1921);
not gate_1818(G580,G1916);
and gate_1819(G1256,G1209,G1231);
and gate_1820(G1261,G1216,G1231);
and gate_1821(G1266,G1223,G1231);
and gate_1822(G1271,G1080,G1231);
not gate_1823(G1486,G1483);
and gate_1824(G1934,G1887,G1909);
and gate_1825(G1942,G1894,G1909);
and gate_1826(G1947,G1901,G1909);
and gate_1827(G1952,G1758,G1909);
not gate_1828(G2163,G2160);
not gate_1829(G5250,G5244);
nand gate_1830(G3537,G5244,G5251);
not gate_1831(G5258,G5252);
nand gate_1832(G3542,G5252,G5259);
and gate_1833(G3782,G1253,G3737,G3765);
and gate_1834(G3785,G1248,G3737,G3765);
and gate_1835(G3788,G1243,G3737,G3765);
or gate_1836(G3790,G3778,G3779,G3780);
and gate_1837(G3843,G1926,G3795,G3823);
and gate_1838(G3846,G1921,G3795,G3823);
or gate_1839(G3849,G3839,G3840,G3841);
nand gate_1840(G3960,G5409,G5412);
not gate_1841(G5413,G5409);
nand gate_1842(G3963,G5417,G5420);
and gate_1843(G4010,G1238,G3972,G3998);
and gate_1844(G4068,G1916,G4030,G4056);
nand gate_1845(G4358,G4356,G4357);
nand gate_1846(G4416,G4414,G4415);
not gate_1847(G4480,G4474);
nand gate_1848(G4483,G4474,G4481);
not gate_1849(G4568,G4562);
nand gate_1850(G4571,G4562,G4569);
nand gate_1851(G4822,G4820,G4821);
nand gate_1852(G4880,G4878,G4879);
nand gate_1853(G4938,G4936,G4937);
not gate_1854(G5022,G5016);
nand gate_1855(G5025,G5016,G5023);
or gate_1856(G1258,G1256,G1257);
or gate_1857(G1263,G1261,G1262);
or gate_1858(G1268,G1266,G1267);
or gate_1859(G1273,G1271,G1272);
or gate_1860(G1936,G1934,G1935);
or gate_1861(G1944,G1942,G1943);
or gate_1862(G1949,G1947,G1948);
or gate_1863(G1954,G1952,G1953);
nand gate_1864(G3536,G5247,G5250);
nand gate_1865(G3541,G5255,G5258);
or gate_1866(G3791,G3781,G3782,G3783);
or gate_1867(G3792,G3784,G3785,G3786);
or gate_1868(G3793,G3787,G3788,G3789);
or gate_1869(G3850,G3842,G3843,G3844);
or gate_1870(G3851,G3845,G3846,G3847);
nand gate_1871(G3961,G5406,G5413);
nand gate_1872(G3965,G3963,G3964);
or gate_1873(G4024,G4009,G4010,G4011);
or gate_1874(G4082,G4067,G4068,G4069);
nand gate_1875(G4482,G4477,G4480);
nand gate_1876(G4570,G4565,G4568);
nand gate_1877(G5024,G5019,G5022);
and gate_1878(G1666,G3790,G1609,G1645);
and gate_1879(G1670,G3849,G1621,G1645);
and gate_1880(G2337,G3790,G2281,G2316);
and gate_1881(G2341,G3849,G2293,G2316);
and gate_1882(G719,G3790,G2418,G2454);
and gate_1883(G758,G3849,G2430,G2454);
and gate_1884(G798,G3849,G2488,G2512);
not gate_1885(G838,G3849);
and gate_1886(G856,G3790,G2476,G2512);
not gate_1887(G861,G3790);
nand gate_1888(G3538,G3536,G3537);
nand gate_1889(G3543,G3541,G3542);
nand gate_1890(G3962,G3960,G3961);
not gate_1891(G4364,G4358);
nand gate_1892(G4367,G4358,G4365);
not gate_1893(G4422,G4416);
nand gate_1894(G4425,G4416,G4423);
nand gate_1895(G4484,G4482,G4483);
nand gate_1896(G4572,G4570,G4571);
not gate_1897(G4828,G4822);
nand gate_1898(G4831,G4822,G4829);
not gate_1899(G4886,G4880);
nand gate_1900(G4889,G4880,G4887);
not gate_1901(G4944,G4938);
nand gate_1902(G4947,G4938,G4945);
nand gate_1903(G5026,G5024,G5025);
not gate_1904(G571,G1273);
not gate_1905(G572,G1268);
not gate_1906(G573,G1263);
not gate_1907(G574,G1258);
not gate_1908(G581,G1954);
not gate_1909(G582,G1949);
not gate_1910(G583,G1944);
not gate_1911(G584,G1936);
not gate_1912(G623,G1936);
and gate_1913(G1576,G4082,G1540,G1564);
and gate_1914(G1578,G4024,G1528,G1564);
or gate_1915(G659,G1664,G1666,G1667,G1668);
and gate_1916(G1672,G3791,G1609,G1645);
and gate_1917(G1676,G3850,G1621,G1645);
and gate_1918(G1678,G3792,G1609,G1645);
and gate_1919(G1682,G3851,G1621,G1645);
and gate_1920(G1684,G3793,G1609,G1645);
and gate_1921(G2250,G4082,G2215,G2238);
and gate_1922(G2252,G4024,G2203,G2238);
or gate_1923(G691,G2335,G2337,G2338,G2339);
and gate_1924(G2343,G3791,G2281,G2316);
and gate_1925(G2347,G3850,G2293,G2316);
and gate_1926(G2349,G3792,G2281,G2316);
and gate_1927(G2353,G3851,G2293,G2316);
and gate_1928(G2355,G3793,G2281,G2316);
or gate_1929(G722,G718,G719,G720,G721);
and gate_1930(G743,G4082,G3570,G3594);
and gate_1931(G744,G4024,G3558,G3594);
and gate_1932(G748,G3851,G2430,G2454);
and gate_1933(G749,G3793,G2418,G2454);
and gate_1934(G753,G3850,G2430,G2454);
and gate_1935(G754,G3792,G2418,G2454);
and gate_1936(G759,G3791,G2418,G2454);
and gate_1937(G783,G4082,G3672,G3696);
and gate_1938(G784,G4024,G3660,G3696);
and gate_1939(G788,G3851,G2488,G2512);
and gate_1940(G789,G3793,G2476,G2512);
and gate_1941(G793,G3850,G2488,G2512);
and gate_1942(G794,G3792,G2476,G2512);
and gate_1943(G799,G3791,G2476,G2512);
and gate_1944(G3735,G1936,G3724,G3717);
not gate_1945(G832,G4082);
not gate_1946(G834,G3851);
not gate_1947(G836,G3850);
not gate_1948(G3835,G3965);
or gate_1949(G859,G855,G856,G857,G858);
not gate_1950(G871,G4024);
not gate_1951(G873,G3793);
not gate_1952(G875,G3792);
not gate_1953(G877,G3791);
buf gate_1954(G998,G3538);
buf gate_1955(G1000,G3543);
and gate_1956(G3651,G3965,G3632);
and gate_1957(G4013,G1273,G3972,G3998);
and gate_1958(G4016,G1268,G3972,G3998);
and gate_1959(G4019,G1263,G3972,G3998);
and gate_1960(G4022,G1258,G3972,G3998);
and gate_1961(G4071,G1954,G4030,G4056);
and gate_1962(G4074,G1949,G4030,G4056);
and gate_1963(G4077,G1944,G4030,G4056);
and gate_1964(G4080,G1936,G4030,G4056);
nand gate_1965(G4096,G4113,G1936);
nand gate_1966(G4366,G4361,G4364);
nand gate_1967(G4424,G4419,G4422);
nand gate_1968(G4830,G4825,G4828);
nand gate_1969(G4888,G4883,G4886);
nand gate_1970(G4946,G4941,G4944);
and gate_1971(G575,G566,G567,G568,G569,G570,G571,G572,G573,G574);
and gate_1972(G585,G576,G577,G578,G579,G580,G581,G582,G583,G584);
or gate_1973(G640,G1576,G1578,G1579,G1580);
and gate_1974(G661,G659,G1606);
or gate_1975(G662,G1670,G1672,G1673,G1674);
or gate_1976(G665,G1676,G1678,G1679,G1680);
or gate_1977(G668,G1682,G1684,G1685,G1686);
or gate_1978(G674,G2250,G2252,G2253,G2254);
and gate_1979(G693,G691,G2279);
or gate_1980(G694,G2341,G2343,G2344,G2345);
or gate_1981(G697,G2347,G2349,G2350,G2351);
or gate_1982(G700,G2353,G2355,G2356,G2357);
or gate_1983(G747,G743,G744,G745,G746);
or gate_1984(G752,G748,G749,G750,G751);
or gate_1985(G757,G753,G754,G755,G756);
or gate_1986(G762,G758,G759,G760,G761);
or gate_1987(G787,G783,G784,G785,G786);
or gate_1988(G792,G788,G789,G790,G791);
or gate_1989(G797,G793,G794,G795,G796);
or gate_1990(G802,G798,G799,G800,G801);
or gate_1991(G817,G3731,G3733,G3734,G3735);
and gate_1992(G839,G3835,G3803,G3823);
not gate_1993(G3540,G3538);
not gate_1994(G3545,G3543);
not gate_1995(G3777,G3962);
and gate_1996(G3648,G3962,G3632);
or gate_1997(G4025,G4012,G4013,G4014);
or gate_1998(G4026,G4015,G4016,G4017);
or gate_1999(G4027,G4018,G4019,G4020);
or gate_2000(G4028,G4021,G4022,G4023);
or gate_2001(G4083,G4070,G4071,G4072);
or gate_2002(G4084,G4073,G4074,G4075);
or gate_2003(G4085,G4076,G4077,G4078);
or gate_2004(G4086,G4079,G4080,G4081);
nand gate_2005(G4368,G4366,G4367);
nand gate_2006(G4426,G4424,G4425);
not gate_2007(G4490,G4484);
nand gate_2008(G4493,G4484,G4491);
not gate_2009(G4578,G4572);
nand gate_2010(G4581,G4572,G4579);
nand gate_2011(G4832,G4830,G4831);
nand gate_2012(G4890,G4888,G4889);
nand gate_2013(G4948,G4946,G4947);
not gate_2014(G5032,G5026);
nand gate_2015(G5035,G5026,G5033);
and gate_2016(G642,G640,G1526);
and gate_2017(G664,G662,G1606);
and gate_2018(G667,G665,G1606);
and gate_2019(G670,G668,G1606);
and gate_2020(G676,G674,G2202);
and gate_2021(G696,G694,G2279);
and gate_2022(G699,G697,G2279);
and gate_2023(G702,G700,G2279);
and gate_2024(G811,G4113,G4096);
and gate_2025(G812,G4096,G1936);
and gate_2026(G818,G816,G817);
and gate_2027(G853,G562,G3540,G3545,G3535,G3970);
and gate_2028(G878,G3777,G3745,G3765);
nand gate_2029(G4492,G4487,G4490);
nand gate_2030(G4580,G4575,G4578);
nand gate_2031(G5034,G5029,G5032);
and gate_2032(G1582,G4083,G1540,G1564);
and gate_2033(G1584,G4025,G1528,G1564);
and gate_2034(G1588,G4084,G1540,G1564);
and gate_2035(G1590,G4026,G1528,G1564);
and gate_2036(G1594,G4085,G1540,G1564);
and gate_2037(G1596,G4027,G1528,G1564);
and gate_2038(G1600,G4086,G1540,G1564);
and gate_2039(G1602,G4028,G1528,G1564);
and gate_2040(G2256,G4083,G2215,G2238);
and gate_2041(G2258,G4025,G2203,G2238);
and gate_2042(G2262,G4084,G2215,G2238);
and gate_2043(G2264,G4026,G2203,G2238);
and gate_2044(G2268,G4085,G2215,G2238);
and gate_2045(G2270,G4027,G2203,G2238);
and gate_2046(G2274,G4086,G2215,G2238);
and gate_2047(G2276,G4028,G2203,G2238);
and gate_2048(G708,G4086,G3672,G3696);
and gate_2049(G709,G4028,G3660,G3696);
and gate_2050(G723,G4086,G3570,G3594);
and gate_2051(G724,G4028,G3558,G3594);
and gate_2052(G728,G4085,G3570,G3594);
and gate_2053(G729,G4027,G3558,G3594);
and gate_2054(G733,G4084,G3570,G3594);
and gate_2055(G734,G4026,G3558,G3594);
and gate_2056(G738,G4083,G3570,G3594);
and gate_2057(G739,G4025,G3558,G3594);
and gate_2058(G768,G4085,G3672,G3696);
and gate_2059(G769,G4027,G3660,G3696);
and gate_2060(G773,G4084,G3672,G3696);
and gate_2061(G774,G4026,G3660,G3696);
and gate_2062(G778,G4083,G3672,G3696);
and gate_2063(G779,G4025,G3660,G3696);
or gate_2064(G813,G811,G812);
not gate_2065(G824,G4086);
not gate_2066(G826,G4085);
not gate_2067(G828,G4084);
not gate_2068(G830,G4083);
and gate_2069(G854,G852,G853,G245);
not gate_2070(G863,G4028);
not gate_2071(G865,G4027);
not gate_2072(G867,G4026);
not gate_2073(G869,G4025);
not gate_2074(G4374,G4368);
nand gate_2075(G4377,G4368,G4375);
not gate_2076(G4432,G4426);
nand gate_2077(G4435,G4426,G4433);
nand gate_2078(G4494,G4492,G4493);
nand gate_2079(G4582,G4580,G4581);
not gate_2080(G4838,G4832);
nand gate_2081(G4841,G4832,G4839);
not gate_2082(G4896,G4890);
nand gate_2083(G4899,G4890,G4897);
not gate_2084(G4954,G4948);
nand gate_2085(G4957,G4948,G4955);
nand gate_2086(G5036,G5034,G5035);
or gate_2087(G643,G1582,G1584,G1585,G1586);
or gate_2088(G646,G1588,G1590,G1591,G1592);
or gate_2089(G649,G1594,G1596,G1597,G1598);
or gate_2090(G652,G1600,G1602,G1603,G1604);
or gate_2091(G677,G2256,G2258,G2259,G2260);
or gate_2092(G680,G2262,G2264,G2265,G2266);
or gate_2093(G683,G2268,G2270,G2271,G2272);
or gate_2094(G686,G2274,G2276,G2277,G2278);
or gate_2095(G712,G708,G709,G710,G711);
or gate_2096(G727,G723,G724,G725,G726);
or gate_2097(G732,G728,G729,G730,G731);
or gate_2098(G737,G733,G734,G735,G736);
or gate_2099(G742,G738,G739,G740,G741);
or gate_2100(G772,G768,G769,G770,G771);
or gate_2101(G777,G773,G774,G775,G776);
or gate_2102(G782,G778,G779,G780,G781);
nand gate_2103(G4376,G4371,G4374);
nand gate_2104(G4434,G4429,G4432);
nand gate_2105(G4840,G4835,G4838);
nand gate_2106(G4898,G4893,G4896);
nand gate_2107(G4956,G4951,G4954);
and gate_2108(G645,G643,G1526);
and gate_2109(G648,G646,G1526);
and gate_2110(G651,G649,G1526);
and gate_2111(G654,G652,G1526);
and gate_2112(G679,G677,G2202);
and gate_2113(G682,G680,G2202);
and gate_2114(G685,G683,G2202);
and gate_2115(G688,G686,G2202);
nand gate_2116(G4378,G4376,G4377);
nand gate_2117(G4436,G4434,G4435);
not gate_2118(G4500,G4494);
nand gate_2119(G4503,G4494,G4501);
not gate_2120(G4588,G4582);
nand gate_2121(G4591,G4582,G4589);
nand gate_2122(G4842,G4840,G4841);
nand gate_2123(G4900,G4898,G4899);
nand gate_2124(G4958,G4956,G4957);
not gate_2125(G5042,G5036);
nand gate_2126(G5045,G5036,G5043);
nand gate_2127(G4502,G4497,G4500);
nand gate_2128(G4590,G4585,G4588);
nand gate_2129(G5044,G5039,G5042);
not gate_2130(G4384,G4378);
nand gate_2131(G4387,G4378,G4385);
not gate_2132(G4442,G4436);
nand gate_2133(G4445,G4436,G4443);
nand gate_2134(G4504,G4502,G4503);
nand gate_2135(G4592,G4590,G4591);
not gate_2136(G4848,G4842);
nand gate_2137(G4851,G4842,G4849);
not gate_2138(G4906,G4900);
nand gate_2139(G4909,G4900,G4907);
not gate_2140(G4964,G4958);
nand gate_2141(G4967,G4958,G4965);
nand gate_2142(G5046,G5044,G5045);
nand gate_2143(G4386,G4381,G4384);
nand gate_2144(G4444,G4439,G4442);
nand gate_2145(G4850,G4845,G4848);
nand gate_2146(G4908,G4903,G4906);
nand gate_2147(G4966,G4961,G4964);
nand gate_2148(G4388,G4386,G4387);
nand gate_2149(G4446,G4444,G4445);
not gate_2150(G4510,G4504);
nand gate_2151(G4513,G4504,G4511);
not gate_2152(G4598,G4592);
nand gate_2153(G4601,G4592,G4599);
nand gate_2154(G4852,G4850,G4851);
nand gate_2155(G4910,G4908,G4909);
nand gate_2156(G4968,G4966,G4967);
not gate_2157(G5052,G5046);
nand gate_2158(G5055,G5046,G5053);
nand gate_2159(G4512,G4507,G4510);
nand gate_2160(G4600,G4595,G4598);
nand gate_2161(G5054,G5049,G5052);
not gate_2162(G4394,G4388);
nand gate_2163(G4397,G4388,G4395);
not gate_2164(G4452,G4446);
nand gate_2165(G4455,G4446,G4453);
nand gate_2166(G4514,G4512,G4513);
nand gate_2167(G4602,G4600,G4601);
not gate_2168(G4858,G4852);
nand gate_2169(G4861,G4852,G4859);
not gate_2170(G4916,G4910);
nand gate_2171(G4919,G4910,G4917);
not gate_2172(G4974,G4968);
nand gate_2173(G4977,G4968,G4975);
nand gate_2174(G5056,G5054,G5055);
nand gate_2175(G4396,G4391,G4394);
nand gate_2176(G4454,G4449,G4452);
nand gate_2177(G4860,G4855,G4858);
nand gate_2178(G4918,G4913,G4916);
nand gate_2179(G4976,G4971,G4974);
nand gate_2180(G4398,G4396,G4397);
nand gate_2181(G4456,G4454,G4455);
not gate_2182(G4520,G4514);
nand gate_2183(G4523,G4514,G4521);
not gate_2184(G4608,G4602);
nand gate_2185(G4611,G4602,G4609);
nand gate_2186(G4862,G4860,G4861);
nand gate_2187(G4920,G4918,G4919);
nand gate_2188(G4978,G4976,G4977);
not gate_2189(G5062,G5056);
nand gate_2190(G5065,G5056,G5063);
nand gate_2191(G4522,G4517,G4520);
nand gate_2192(G4610,G4605,G4608);
nand gate_2193(G5064,G5059,G5062);
not gate_2194(G4404,G4398);
nand gate_2195(G1488,G4398,G4405);
not gate_2196(G4462,G4456);
nand gate_2197(G1493,G4456,G4463);
not gate_2198(G4868,G4862);
nand gate_2199(G2165,G4862,G4869);
not gate_2200(G4926,G4920);
nand gate_2201(G2170,G4920,G4927);
nand gate_2202(G4524,G4522,G4523);
nand gate_2203(G4612,G4610,G4611);
not gate_2204(G4984,G4978);
nand gate_2205(G4987,G4978,G4985);
nand gate_2206(G5066,G5064,G5065);
nand gate_2207(G1487,G4401,G4404);
nand gate_2208(G1492,G4459,G4462);
nand gate_2209(G2164,G4865,G4868);
nand gate_2210(G2169,G4923,G4926);
nand gate_2211(G4986,G4981,G4984);
nand gate_2212(G1489,G1487,G1488);
nand gate_2213(G1494,G1492,G1493);
nand gate_2214(G2166,G2164,G2165);
nand gate_2215(G2171,G2169,G2170);
not gate_2216(G4530,G4524);
nand gate_2217(G4533,G4524,G4531);
not gate_2218(G4618,G4612);
nand gate_2219(G4543,G4612,G4619);
nand gate_2220(G4988,G4986,G4987);
not gate_2221(G5072,G5066);
nand gate_2222(G4997,G5066,G5073);
nand gate_2223(G4532,G4527,G4530);
nand gate_2224(G4542,G4615,G4618);
nand gate_2225(G4996,G5069,G5072);
and gate_2226(G1513,G1494,G1462,G1502);
and gate_2227(G1514,G1489,G1458,G1502);
and gate_2228(G1515,G1494,G1483,G1497);
and gate_2229(G1516,G1489,G1486,G1497);
not gate_2230(G4994,G4988);
nand gate_2231(G2184,G4988,G4995);
and gate_2232(G2190,G2171,G2139,G2179);
and gate_2233(G2191,G2166,G2135,G2179);
and gate_2234(G2192,G2171,G2160,G2174);
and gate_2235(G2193,G2166,G2163,G2174);
nand gate_2236(G4534,G4532,G4533);
nand gate_2237(G4544,G4542,G4543);
nand gate_2238(G4998,G4996,G4997);
nand gate_2239(G2183,G4991,G4994);
or gate_2240(G4620,G1513,G1514,G1515,G1516);
or gate_2241(G5074,G2190,G2191,G2192,G2193);
not gate_2242(G4540,G4534);
nand gate_2243(G1507,G4534,G4541);
not gate_2244(G4550,G4544);
nand gate_2245(G1510,G4544,G4551);
nand gate_2246(G2185,G2183,G2184);
not gate_2247(G5004,G4998);
nand gate_2248(G2187,G4998,G5005);
nand gate_2249(G1506,G4537,G4540);
nand gate_2250(G1509,G4547,G4550);
not gate_2251(G4626,G4620);
nand gate_2252(G2186,G5001,G5004);
and gate_2253(G2195,G2174,G2185);
not gate_2254(G5080,G5074);
nand gate_2255(G1508,G1506,G1507);
nand gate_2256(G1511,G1509,G1510);
nand gate_2257(G2188,G2186,G2187);
not gate_2258(G1512,G1511);
and gate_2259(G1518,G1497,G1508);
not gate_2260(G2189,G2188);
and gate_2261(G1517,G1512,G1502);
and gate_2262(G2194,G2189,G2179);
or gate_2263(G4623,G1517,G1518);
or gate_2264(G5077,G2194,G2195);
nand gate_2265(G1519,G4623,G4626);
not gate_2266(G4627,G4623);
nand gate_2267(G2196,G5077,G5080);
not gate_2268(G5081,G5077);
nand gate_2269(G1520,G4620,G4627);
nand gate_2270(G2197,G5074,G5081);
nand gate_2271(G1521,G1519,G1520);
nand gate_2272(G2198,G2196,G2197);
and gate_2273(G840,G2198,G3795,G3823);
and gate_2274(G879,G1521,G3737,G3765);
not gate_2275(G1524,G1521);
not gate_2276(G2201,G2198);
or gate_2277(G843,G839,G840,G841,G842);
or gate_2278(G882,G878,G879,G880,G881);
and gate_2279(G3649,G1524,G3628);
and gate_2280(G3652,G2201,G3628);
or gate_2281(G3657,G3648,G3649);
or gate_2282(G3658,G3651,G3652);
and gate_2283(G3636,G3657,G3622);
and gate_2284(G3639,G3658,G3622);
and gate_2285(G3642,G3657,G3622);
and gate_2286(G3645,G3658,G3622);
or gate_2287(G3653,G3636,G3637);
or gate_2288(G3654,G3639,G3640);
or gate_2289(G3655,G3642,G3643);
or gate_2290(G3656,G3645,G3646);
and gate_2291(G763,G3656,G2430,G2454);
and gate_2292(G764,G3655,G2418,G2454);
and gate_2293(G803,G3656,G2488,G2512);
and gate_2294(G804,G3655,G2476,G2512);
and gate_2295(G1657,G3654,G1621,G1645);
and gate_2296(G1659,G3653,G1609,G1645);
and gate_2297(G2328,G3654,G2293,G2316);
and gate_2298(G2330,G3653,G2281,G2316);
or gate_2299(G1662,G1657,G1659,G1660,G1661);
or gate_2300(G2333,G2328,G2330,G2331,G2332);
or gate_2301(G767,G763,G764,G765,G766);
or gate_2302(G807,G803,G804,G805,G806);
and gate_2303(G657,G1662,G1606);
and gate_2304(G689,G2333,G2279);
not gate_2305(G658,G657);
not gate_2306(G690,G689);
endmodule
