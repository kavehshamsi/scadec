// Verilog File 
module i4 (pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,pi133,pi134,pi135,pi136,pi137,pi138,
pi139,pi140,pi141,pi142,pi143,pi144,pi145,pi146,pi147,pi148,
pi149,pi150,pi151,pi152,pi153,pi154,pi155,pi156,pi157,pi158,
pi159,pi160,pi161,pi162,pi163,pi164,pi165,pi166,pi167,pi168,
pi169,pi170,pi171,pi172,pi173,pi174,pi175,pi176,pi177,pi178,
pi179,pi180,pi181,pi182,pi183,pi184,pi185,pi186,pi187,pi188,
pi189,pi190,pi191,po0,po1,po2,po3,po4,po5);

input pi000,pi001,pi002,pi003,pi004,pi005,pi006,pi007,pi008,
pi009,pi010,pi011,pi012,pi013,pi014,pi015,pi016,pi017,pi018,
pi019,pi020,pi021,pi022,pi023,pi024,pi025,pi026,pi027,pi028,
pi029,pi030,pi031,pi032,pi033,pi034,pi035,pi036,pi037,pi038,
pi039,pi040,pi041,pi042,pi043,pi044,pi045,pi046,pi047,pi048,
pi049,pi050,pi051,pi052,pi053,pi054,pi055,pi056,pi057,pi058,
pi059,pi060,pi061,pi062,pi063,pi064,pi065,pi066,pi067,pi068,
pi069,pi070,pi071,pi072,pi073,pi074,pi075,pi076,pi077,pi078,
pi079,pi080,pi081,pi082,pi083,pi084,pi085,pi086,pi087,pi088,
pi089,pi090,pi091,pi092,pi093,pi094,pi095,pi096,pi097,pi098,
pi099,pi100,pi101,pi102,pi103,pi104,pi105,pi106,pi107,pi108,
pi109,pi110,pi111,pi112,pi113,pi114,pi115,pi116,pi117,pi118,
pi119,pi120,pi121,pi122,pi123,pi124,pi125,pi126,pi127,pi128,
pi129,pi130,pi131,pi132,pi133,pi134,pi135,pi136,pi137,pi138,
pi139,pi140,pi141,pi142,pi143,pi144,pi145,pi146,pi147,pi148,
pi149,pi150,pi151,pi152,pi153,pi154,pi155,pi156,pi157,pi158,
pi159,pi160,pi161,pi162,pi163,pi164,pi165,pi166,pi167,pi168,
pi169,pi170,pi171,pi172,pi173,pi174,pi175,pi176,pi177,pi178,
pi179,pi180,pi181,pi182,pi183,pi184,pi185,pi186,pi187,pi188,
pi189,pi190,pi191;

output po0,po1,po2,po3,po4,po5;

wire n200,n201,n202,n203,n204,n205,n206,n207,n208,
n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,
n219,n220,n221,n222,n223,n224,n225,n226,n227,n228,
n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,
n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,
n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,
n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,
n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,
n279,n280,n281,n282,n284,n285,n286,n287,n288,n289,
n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,
n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,
n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,
n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,
n330,n331,n332,n333,n334,n335,n336,n337,n338,n339,
n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,
n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,
n360,n361,n362,n363,n364,n365,n366,n368,n369,n370,
n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,
n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,
n391,n392,n393,n394,n395,n396,n397,n398,n399,n400,
n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,
n411,n412,n413,n414,n415,n416,n417,n418,n419,n420,
n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,
n431,n432,n433,n434,n435,n436,n437,n438,n439,n440,
n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,
n452,n453,n454,n455,n456,n457,n458,n459,n460,n461,
n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,
n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,
n482,n483,n484,n485,n486,n487,n488,n489,n490,n491,
n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,
n502,n503,n504,n505,n506,n507,n508,n509,n510,n511,
n512,n513,n514,n515,n516,n517,n518,n519,n520,n521,
n522,n523,n524,n525,n526,n527,n528,n529,n530,n531,
n532,n533,n534;
and gate_0(po0,pi000,pi001);
and gate_1(po1,pi002,pi003);
and gate_2(n200,pi039,pi040);
and gate_3(n201,pi041,n200);
and gate_4(n202,pi036,n201);
not gate_5(n203,n202);
and gate_6(n204,pi004,pi005);
not gate_7(n205,n204);
and gate_8(n206,n203,n205);
and gate_9(n207,pi010,pi011);
not gate_10(n208,n207);
and gate_11(n209,pi066,pi067);
and gate_12(n210,pi068,n209);
and gate_13(n211,pi063,n210);
not gate_14(n212,n211);
and gate_15(n213,n208,n212);
and gate_16(n214,pi063,pi069);
and gate_17(n215,pi070,n214);
and gate_18(n216,pi071,n215);
and gate_19(n217,pi066,n216);
not gate_20(n218,n217);
and gate_21(n219,pi063,pi064);
and gate_22(n220,pi065,n219);
not gate_23(n221,n220);
and gate_24(n222,n218,n221);
and gate_25(n223,n213,n222);
not gate_26(n224,n223);
and gate_27(n225,pi180,pi182);
and gate_28(n226,n224,n225);
and gate_29(n227,pi181,n226);
not gate_30(n228,n227);
and gate_31(n229,pi006,pi007);
not gate_32(n230,n229);
and gate_33(n231,pi048,pi049);
and gate_34(n232,pi050,n231);
and gate_35(n233,pi045,n232);
not gate_36(n234,n233);
and gate_37(n235,n230,n234);
and gate_38(n236,pi045,pi051);
and gate_39(n237,pi052,n236);
and gate_40(n238,pi053,n237);
and gate_41(n239,pi048,n238);
not gate_42(n240,n239);
and gate_43(n241,pi045,pi046);
and gate_44(n242,pi047,n241);
not gate_45(n243,n242);
and gate_46(n244,n240,n243);
and gate_47(n245,n235,n244);
not gate_48(n246,n245);
and gate_49(n247,pi180,n246);
not gate_50(n248,n247);
and gate_51(n249,n228,n248);
and gate_52(n250,n206,n249);
and gate_53(n251,pi008,pi009);
not gate_54(n252,n251);
and gate_55(n253,pi057,pi058);
and gate_56(n254,pi059,n253);
and gate_57(n255,pi054,n254);
not gate_58(n256,n255);
and gate_59(n257,n252,n256);
and gate_60(n258,pi054,pi060);
and gate_61(n259,pi061,n258);
and gate_62(n260,pi062,n259);
and gate_63(n261,pi057,n260);
not gate_64(n262,n261);
and gate_65(n263,pi054,pi055);
and gate_66(n264,pi056,n263);
not gate_67(n265,n264);
and gate_68(n266,n262,n265);
and gate_69(n267,n257,n266);
not gate_70(n268,n267);
and gate_71(n269,pi181,n268);
and gate_72(n270,pi180,n269);
not gate_73(n271,n270);
and gate_74(n272,pi036,pi037);
and gate_75(n273,pi038,n272);
not gate_76(n274,n273);
and gate_77(n275,pi036,pi042);
and gate_78(n276,pi043,n275);
and gate_79(n277,pi044,n276);
and gate_80(n278,pi039,n277);
not gate_81(n279,n278);
and gate_82(n280,n274,n279);
and gate_83(n281,n271,n280);
and gate_84(n282,n250,n281);
not gate_85(po2,n282);
and gate_86(n284,pi075,pi076);
and gate_87(n285,pi077,n284);
and gate_88(n286,pi072,n285);
not gate_89(n287,n286);
and gate_90(n288,pi012,pi013);
not gate_91(n289,n288);
and gate_92(n290,n287,n289);
and gate_93(n291,pi018,pi019);
not gate_94(n292,n291);
and gate_95(n293,pi102,pi103);
and gate_96(n294,pi104,n293);
and gate_97(n295,pi099,n294);
not gate_98(n296,n295);
and gate_99(n297,n292,n296);
and gate_100(n298,pi099,pi105);
and gate_101(n299,pi106,n298);
and gate_102(n300,pi107,n299);
and gate_103(n301,pi102,n300);
not gate_104(n302,n301);
and gate_105(n303,pi099,pi100);
and gate_106(n304,pi101,n303);
not gate_107(n305,n304);
and gate_108(n306,n302,n305);
and gate_109(n307,n297,n306);
not gate_110(n308,n307);
and gate_111(n309,pi183,pi185);
and gate_112(n310,n308,n309);
and gate_113(n311,pi184,n310);
not gate_114(n312,n311);
and gate_115(n313,pi014,pi015);
not gate_116(n314,n313);
and gate_117(n315,pi084,pi085);
and gate_118(n316,pi086,n315);
and gate_119(n317,pi081,n316);
not gate_120(n318,n317);
and gate_121(n319,n314,n318);
and gate_122(n320,pi081,pi087);
and gate_123(n321,pi088,n320);
and gate_124(n322,pi089,n321);
and gate_125(n323,pi084,n322);
not gate_126(n324,n323);
and gate_127(n325,pi081,pi082);
and gate_128(n326,pi083,n325);
not gate_129(n327,n326);
and gate_130(n328,n324,n327);
and gate_131(n329,n319,n328);
not gate_132(n330,n329);
and gate_133(n331,pi183,n330);
not gate_134(n332,n331);
and gate_135(n333,n312,n332);
and gate_136(n334,n290,n333);
and gate_137(n335,pi016,pi017);
not gate_138(n336,n335);
and gate_139(n337,pi093,pi094);
and gate_140(n338,pi095,n337);
and gate_141(n339,pi090,n338);
not gate_142(n340,n339);
and gate_143(n341,n336,n340);
and gate_144(n342,pi090,pi096);
and gate_145(n343,pi097,n342);
and gate_146(n344,pi098,n343);
and gate_147(n345,pi093,n344);
not gate_148(n346,n345);
and gate_149(n347,pi090,pi091);
and gate_150(n348,pi092,n347);
not gate_151(n349,n348);
and gate_152(n350,n346,n349);
and gate_153(n351,n341,n350);
not gate_154(n352,n351);
and gate_155(n353,pi184,n352);
and gate_156(n354,pi183,n353);
not gate_157(n355,n354);
and gate_158(n356,pi072,pi073);
and gate_159(n357,pi074,n356);
not gate_160(n358,n357);
and gate_161(n359,pi072,pi078);
and gate_162(n360,pi079,n359);
and gate_163(n361,pi080,n360);
and gate_164(n362,pi075,n361);
not gate_165(n363,n362);
and gate_166(n364,n358,n363);
and gate_167(n365,n355,n364);
and gate_168(n366,n334,n365);
not gate_169(po3,n366);
and gate_170(n368,pi111,pi112);
and gate_171(n369,pi113,n368);
and gate_172(n370,pi108,n369);
not gate_173(n371,n370);
and gate_174(n372,pi020,pi021);
not gate_175(n373,n372);
and gate_176(n374,n371,n373);
and gate_177(n375,pi026,pi027);
not gate_178(n376,n375);
and gate_179(n377,pi138,pi139);
and gate_180(n378,pi140,n377);
and gate_181(n379,pi135,n378);
not gate_182(n380,n379);
and gate_183(n381,n376,n380);
and gate_184(n382,pi135,pi141);
and gate_185(n383,pi142,n382);
and gate_186(n384,pi143,n383);
and gate_187(n385,pi138,n384);
not gate_188(n386,n385);
and gate_189(n387,pi135,pi136);
and gate_190(n388,pi137,n387);
not gate_191(n389,n388);
and gate_192(n390,n386,n389);
and gate_193(n391,n381,n390);
not gate_194(n392,n391);
and gate_195(n393,pi186,pi188);
and gate_196(n394,n392,n393);
and gate_197(n395,pi187,n394);
not gate_198(n396,n395);
and gate_199(n397,pi022,pi023);
not gate_200(n398,n397);
and gate_201(n399,pi120,pi121);
and gate_202(n400,pi122,n399);
and gate_203(n401,pi117,n400);
not gate_204(n402,n401);
and gate_205(n403,n398,n402);
and gate_206(n404,pi117,pi123);
and gate_207(n405,pi124,n404);
and gate_208(n406,pi125,n405);
and gate_209(n407,pi120,n406);
not gate_210(n408,n407);
and gate_211(n409,pi117,pi118);
and gate_212(n410,pi119,n409);
not gate_213(n411,n410);
and gate_214(n412,n408,n411);
and gate_215(n413,n403,n412);
not gate_216(n414,n413);
and gate_217(n415,pi186,n414);
not gate_218(n416,n415);
and gate_219(n417,n396,n416);
and gate_220(n418,n374,n417);
and gate_221(n419,pi024,pi025);
not gate_222(n420,n419);
and gate_223(n421,pi129,pi130);
and gate_224(n422,pi131,n421);
and gate_225(n423,pi126,n422);
not gate_226(n424,n423);
and gate_227(n425,n420,n424);
and gate_228(n426,pi126,pi132);
and gate_229(n427,pi133,n426);
and gate_230(n428,pi134,n427);
and gate_231(n429,pi129,n428);
not gate_232(n430,n429);
and gate_233(n431,pi126,pi127);
and gate_234(n432,pi128,n431);
not gate_235(n433,n432);
and gate_236(n434,n430,n433);
and gate_237(n435,n425,n434);
not gate_238(n436,n435);
and gate_239(n437,pi187,n436);
and gate_240(n438,pi186,n437);
not gate_241(n439,n438);
and gate_242(n440,pi108,pi109);
and gate_243(n441,pi110,n440);
not gate_244(n442,n441);
and gate_245(n443,pi108,pi114);
and gate_246(n444,pi115,n443);
and gate_247(n445,pi116,n444);
and gate_248(n446,pi111,n445);
not gate_249(n447,n446);
and gate_250(n448,n442,n447);
and gate_251(n449,n439,n448);
and gate_252(n450,n418,n449);
not gate_253(po4,n450);
and gate_254(n452,pi147,pi148);
and gate_255(n453,pi149,n452);
and gate_256(n454,pi144,n453);
not gate_257(n455,n454);
and gate_258(n456,pi028,pi029);
not gate_259(n457,n456);
and gate_260(n458,n455,n457);
and gate_261(n459,pi034,pi035);
not gate_262(n460,n459);
and gate_263(n461,pi174,pi175);
and gate_264(n462,pi176,n461);
and gate_265(n463,pi171,n462);
not gate_266(n464,n463);
and gate_267(n465,n460,n464);
and gate_268(n466,pi171,pi177);
and gate_269(n467,pi178,n466);
and gate_270(n468,pi179,n467);
and gate_271(n469,pi174,n468);
not gate_272(n470,n469);
and gate_273(n471,pi171,pi172);
and gate_274(n472,pi173,n471);
not gate_275(n473,n472);
and gate_276(n474,n470,n473);
and gate_277(n475,n465,n474);
not gate_278(n476,n475);
and gate_279(n477,pi189,pi191);
and gate_280(n478,n476,n477);
and gate_281(n479,pi190,n478);
not gate_282(n480,n479);
and gate_283(n481,pi030,pi031);
not gate_284(n482,n481);
and gate_285(n483,pi156,pi157);
and gate_286(n484,pi158,n483);
and gate_287(n485,pi153,n484);
not gate_288(n486,n485);
and gate_289(n487,n482,n486);
and gate_290(n488,pi153,pi159);
and gate_291(n489,pi160,n488);
and gate_292(n490,pi161,n489);
and gate_293(n491,pi156,n490);
not gate_294(n492,n491);
and gate_295(n493,pi153,pi154);
and gate_296(n494,pi155,n493);
not gate_297(n495,n494);
and gate_298(n496,n492,n495);
and gate_299(n497,n487,n496);
not gate_300(n498,n497);
and gate_301(n499,pi189,n498);
not gate_302(n500,n499);
and gate_303(n501,n480,n500);
and gate_304(n502,n458,n501);
and gate_305(n503,pi032,pi033);
not gate_306(n504,n503);
and gate_307(n505,pi165,pi166);
and gate_308(n506,pi167,n505);
and gate_309(n507,pi162,n506);
not gate_310(n508,n507);
and gate_311(n509,n504,n508);
and gate_312(n510,pi162,pi168);
and gate_313(n511,pi169,n510);
and gate_314(n512,pi170,n511);
and gate_315(n513,pi165,n512);
not gate_316(n514,n513);
and gate_317(n515,pi162,pi163);
and gate_318(n516,pi164,n515);
not gate_319(n517,n516);
and gate_320(n518,n514,n517);
and gate_321(n519,n509,n518);
not gate_322(n520,n519);
and gate_323(n521,pi190,n520);
and gate_324(n522,pi189,n521);
not gate_325(n523,n522);
and gate_326(n524,pi144,pi145);
and gate_327(n525,pi146,n524);
not gate_328(n526,n525);
and gate_329(n527,pi144,pi150);
and gate_330(n528,pi151,n527);
and gate_331(n529,pi152,n528);
and gate_332(n530,pi147,n529);
not gate_333(n531,n530);
and gate_334(n532,n526,n531);
and gate_335(n533,n523,n532);
and gate_336(n534,n502,n533);
not gate_337(po5,n534);
endmodule
