// Verilog File 
module ex5 (pi0,pi1,pi2,pi3,pi4,pi5,pi6,pi7,po00,
po01,po02,po03,po04,po05,po06,po07,po08,po09,po10,
po11,po12,po13,po14,po15,po16,po17,po18,po19,po20,
po21,po22,po23,po24,po25,po26,po27,po28,po29,po30,
po31,po32,po33,po34,po35,po36,po37,po38,po39,po40,
po41,po42,po43,po44,po45,po46,po47,po48,po49,po50,
po51,po52,po53,po54,po55,po56,po57,po58,po59,po60,
po61,po62);

input pi0,pi1,pi2,pi3,pi4,pi5,pi6,pi7;

output po00,po01,po02,po03,po04,po05,po06,po07,po08,
po09,po10,po11,po12,po13,po14,po15,po16,po17,po18,
po19,po20,po21,po22,po23,po24,po25,po26,po27,po28,
po29,po30,po31,po32,po33,po34,po35,po36,po37,po38,
po39,po40,po41,po42,po43,po44,po45,po46,po47,po48,
po49,po50,po51,po52,po53,po54,po55,po56,po57,po58,
po59,po60,po61,po62;

wire n71,n72,n73,n74,n75,n76,n77,n78,n79,
n80,n82,n83,n85,n86,n87,n88,n89,n92,n93,
n94,n95,n96,n98,n99,n101,n102,n103,n104,n105,
n106,n108,n109,n110,n111,n112,n113,n114,n115,n117,
n118,n119,n120,n121,n122,n123,n124,n125,n126,n128,
n129,n130,n131,n132,n133,n134,n135,n136,n138,n139,
n140,n142,n143,n144,n146,n147,n148,n149,n151,n152,
n153,n155,n156,n158,n159,n160,n162,n163,n165,n166,
n167,n168,n169,n171,n172,n173,n174,n175,n176,n178,
n179,n180,n182,n183,n184,n185,n186,n187,n190,n192,
n193,n194,n196,n197,n199,n201,n202,n203,n204,n206,
n207,n208,n210,n211,n212,n213,n214,n216,n218,n220,
n221,n222,n223,n224,n225,n226,n227,n228,n229,n230,
n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,
n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,
n251,n252,n253,n254,n255,n257,n258,n259,n260,n261,
n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,
n272,n273,n274,n275,n276,n277,n278,n279,n280,n281,
n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,
n292,n293,n294,n295,n296,n298,n299,n300,n301,n302,
n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,
n313,n315,n316,n317,n318,n319,n320,n321,n322,n323,
n324,n325,n326,n327,n328,n329,n330,n331,n332,n333,
n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,
n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,
n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,
n364,n365,n366,n367,n369,n370,n371,n372,n373,n374,
n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,
n386,n387,n388,n389,n390,n391,n392,n393,n394,n395,
n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,
n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,
n417,n418,n419,n420,n421,n422,n423,n424,n425,n426,
n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,
n437,n438,n439,n440,n442,n443,n444,n445,n446,n447,
n448,n449,n450,n451,n452,n453,n454,n455,n456,n457,
n458,n459,n460,n461,n462,n463,n464,n466,n467,n468,
n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,
n479,n480,n481,n482,n483,n484,n485,n486,n487,n488,
n489,n491,n492,n493,n494,n495,n496,n497,n498,n499,
n500,n501,n502,n503,n504,n505,n506,n507,n508,n509,
n510,n511,n512,n513,n514,n515,n516,n517,n518,n519,
n520,n521,n522,n523,n524,n525,n526,n527,n528,n529,
n530,n531,n532,n533,n534,n535,n536,n537,n538,n539,
n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,
n550,n551,n552,n553,n554,n555,n556,n557,n558,n559,
n560,n561,n562,n564,n565,n566,n567,n568,n569,n570,
n571,n572,n573,n574,n575,n576,n578,n579,n580,n581,
n582,n583,n584,n585,n586,n588,n589,n590,n591,n592,
n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,
n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,
n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,
n623,n624,n625,n626,n627,n628,n629,n630,n631,n632,
n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,
n643,n644,n645,n646,n647,n648,n649,n650,n651,n653,
n654,n655,n656,n657,n658,n659,n661,n662,n663,n664,
n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,
n675,n676,n677,n678,n679,n680,n682,n683,n684,n685,
n686,n688,n689,n690,n691,n692,n693,n694,n695,n696,
n697,n698,n699,n700,n701,n702,n703,n704,n705,n706,
n707,n708,n709,n710,n711,n712,n713,n714,n715,n716,
n717,n718,n719,n720,n721,n722,n723,n724,n725,n726,
n727,n729,n730,n731,n732,n733,n735,n736,n737,n738,
n739,n740,n741,n742,n743,n744,n745,n747,n748,n749,
n750,n751,n753,n754,n755,n756,n757,n758,n759,n760,
n761,n762,n763,n764,n765,n766,n767,n768,n769,n770,
n771,n772,n773,n774,n775,n776,n777,n778,n779,n780,
n781,n782,n783,n784,n785,n786,n787,n788,n789,n790,
n791,n792,n793,n795,n796,n797,n798,n799,n800,n801,
n802,n803,n804,n805,n806,n807,n808,n809,n810,n811,
n812,n813,n815,n816,n817,n818,n819,n820,n821,n822,
n823,n824,n825,n826,n827,n828,n829,n830,n831,n832,
n833,n834,n835,n836,n837,n838,n839,n840,n841,n842,
n843,n844,n845,n846,n847,n848,n849,n850,n851,n852,
n853,n854,n855,n856,n857,n858,n859,n860,n861,n862,
n863,n864,n865,n866,n867,n868,n869,n870,n871,n872,
n873,n874,n875,n876,n877,n878,n879,n880,n881,n883,
n884,n885,n886,n887,n888,n889,n890,n891,n892,n893,
n894,n895,n896,n897,n898,n899,n900,n901,n902,n903,
n904,n905,n906,n907,n908,n909,n910,n911,n912,n913,
n914,n915,n916,n917,n918,n919,n920,n921,n922,n923,
n924,n925,n926,n927,n928,n929,n930,n931,n932,n933,
n935,n936,n937,n938,n939,n940,n941,n942,n943,n944,
n945,n946,n947,n948,n949,n950,n951,n952,n953,n954,
n955,n956,n957,n958,n959,n960,n961,n962,n963,n965,
n966,n967,n968,n969,n970,n971,n972,n973,n974,n975,
n976,n977,n978,n979,n980,n981,n982,n983,n984,n985,
n986,n987,n988,n989,n990,n991,n993,n994,n995,n996,
n997,n998,n999,n1000,n1001,n1002,n1003,n1004,n1005,n1006,
n1007,n1008,n1009,n1010,n1011,n1012,n1013,n1014,n1015,n1016,
n1017,n1018,n1019,n1020,n1021,n1022,n1023,n1024,n1025,n1026,
n1027,n1028,n1029,n1030,n1031,n1032,n1033,n1034,n1035,n1036,
n1037,n1038,n1039,n1041,n1042,n1043,n1044,n1045,n1046,n1047,
n1048,n1049,n1050,n1051,n1052,n1053,n1055,n1056,n1057,n1058,
n1059,n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,
n1069,n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,
n1079,n1080,n1081,n1082,n1083,n1084,n1085,n1086,n1087,n1088,
n1089,n1090,n1091,n1092,n1093,n1094,n1095,n1096,n1097,n1098,
n1099,n1100,n1101,n1102,n1104,n1105,n1106,n1107,n1108,n1109,
n1110,n1111,n1112,n1113,n1114,n1115,n1116,n1117,n1119,n1120,
n1121,n1123,n1124;
not gate_0(n71,pi0);
not gate_1(n72,pi1);
not gate_2(n73,pi2);
not gate_3(n74,pi3);
not gate_4(n75,pi4);
not gate_5(n76,pi5);
not gate_6(n77,pi6);
not gate_7(n78,pi7);
and gate_8(n79,n76,n77);
not gate_9(n80,n79);
and gate_10(po00,n75,n79);
not gate_11(n82,po00);
and gate_12(n83,n77,n78);
and gate_13(po01,n76,n83);
and gate_14(n85,pi5,n77);
not gate_15(n86,n85);
and gate_16(n87,n75,n78);
not gate_17(n88,n87);
and gate_18(n89,n85,n87);
and gate_19(po02,n74,n89);
and gate_20(po03,pi3,n89);
and gate_21(n92,pi6,n78);
not gate_22(n93,n92);
and gate_23(n94,n75,n76);
not gate_24(n95,n94);
and gate_25(n96,n92,n94);
and gate_26(po04,pi3,n96);
and gate_27(n98,n75,pi5);
not gate_28(n99,n98);
and gate_29(po05,n92,n98);
not gate_30(n101,po05);
and gate_31(n102,pi3,po00);
not gate_32(n103,n102);
and gate_33(n104,n72,pi2);
not gate_34(n105,n104);
and gate_35(n106,n71,n104);
and gate_36(po06,n102,n106);
and gate_37(n108,n71,pi1);
not gate_38(n109,n108);
and gate_39(n110,n73,n74);
not gate_40(n111,n110);
and gate_41(n112,n108,n110);
and gate_42(n113,n75,n112);
and gate_43(n114,pi6,pi7);
and gate_44(n115,pi5,n114);
and gate_45(po07,n113,n115);
and gate_46(n117,pi1,pi2);
not gate_47(n118,n117);
and gate_48(n119,pi0,n117);
not gate_49(n120,n119);
and gate_50(n121,pi5,pi6);
not gate_51(n122,n121);
and gate_52(n123,n74,n75);
and gate_53(n124,n121,n123);
and gate_54(n125,n119,n124);
not gate_55(n126,n125);
and gate_56(po08,pi7,n125);
and gate_57(n128,n76,n114);
and gate_58(n129,n71,n72);
not gate_59(n130,n129);
and gate_60(n131,pi2,n74);
not gate_61(n132,n131);
and gate_62(n133,n129,n131);
not gate_63(n134,n133);
and gate_64(n135,n75,n133);
not gate_65(n136,n135);
and gate_66(po09,n128,n135);
and gate_67(n138,n98,n114);
and gate_68(n139,n71,n117);
not gate_69(n140,n139);
and gate_70(po10,n138,n139);
and gate_71(n142,pi0,pi1);
not gate_72(n143,n142);
and gate_73(n144,n110,n142);
and gate_74(po11,n138,n144);
and gate_75(n146,pi0,n72);
not gate_76(n147,n146);
and gate_77(n148,n131,n146);
not gate_78(n149,n148);
and gate_79(po12,n138,n148);
and gate_80(n151,n73,pi3);
not gate_81(n152,n151);
and gate_82(n153,n108,n151);
and gate_83(po13,n138,n153);
and gate_84(n155,n146,n151);
not gate_85(n156,n155);
and gate_86(po14,n138,n155);
and gate_87(n158,pi2,n108);
and gate_88(n159,pi3,n98);
and gate_89(n160,n158,n159);
and gate_90(po15,n114,n160);
and gate_91(n162,n142,n151);
not gate_92(n163,n162);
and gate_93(po16,n138,n162);
and gate_94(n165,pi0,n73);
not gate_95(n166,n165);
and gate_96(n167,pi4,n76);
not gate_97(n168,n167);
and gate_98(n169,n72,n167);
and gate_99(po17,n165,n169);
and gate_100(n171,pi2,n76);
not gate_101(n172,n171);
and gate_102(n173,n71,n171);
not gate_103(n174,n173);
and gate_104(n175,pi3,pi4);
and gate_105(n176,n72,n175);
and gate_106(po18,n173,n176);
and gate_107(n178,n74,pi4);
not gate_108(n179,n178);
and gate_109(n180,n73,n178);
and gate_110(po19,n129,n180);
and gate_111(n182,n79,n123);
not gate_112(n183,n182);
and gate_113(n184,n72,n73);
not gate_114(n185,n184);
and gate_115(n186,pi0,n184);
not gate_116(n187,n186);
and gate_117(po20,n182,n186);
and gate_118(po21,n102,n186);
and gate_119(n190,n94,n114);
and gate_120(po22,n186,n190);
not gate_121(n192,po22);
and gate_122(n193,pi3,pi5);
and gate_123(n194,n73,n193);
and gate_124(po23,n129,n194);
and gate_125(n196,n110,n129);
and gate_126(n197,n94,n196);
and gate_127(po24,n92,n197);
and gate_128(n199,n76,n92);
and gate_129(po25,n113,n199);
not gate_130(n201,po25);
and gate_131(n202,pi0,n74);
not gate_132(n203,n202);
and gate_133(n204,pi2,n190);
and gate_134(po26,n202,n204);
and gate_135(n206,n74,n94);
not gate_136(n207,n206);
and gate_137(n208,n158,n206);
and gate_138(po27,n92,n208);
and gate_139(n210,pi3,n75);
not gate_140(n211,n210);
and gate_141(n212,pi2,n210);
not gate_142(n213,n212);
and gate_143(n214,n146,n212);
and gate_144(po28,n128,n214);
and gate_145(n216,n77,pi7);
and gate_146(po29,n197,n216);
and gate_147(n218,n119,n206);
and gate_148(po30,n114,n218);
and gate_149(n220,n99,n168);
not gate_150(n221,n220);
and gate_151(n222,pi4,pi5);
not gate_152(n223,n222);
and gate_153(n224,n95,n223);
not gate_154(n225,n224);
and gate_155(n226,pi0,n104);
not gate_156(n227,n226);
and gate_157(n228,n72,n227);
not gate_158(n229,n228);
and gate_159(n230,n132,n152);
not gate_160(n231,n230);
and gate_161(n232,n129,n231);
not gate_162(n233,n232);
and gate_163(n234,n228,n233);
not gate_164(n235,n234);
and gate_165(n236,n225,n235);
not gate_166(n237,n236);
and gate_167(n238,pi2,pi3);
not gate_168(n239,n238);
and gate_169(n240,n111,n239);
not gate_170(n241,n240);
and gate_171(n242,n72,n241);
not gate_172(n243,n242);
and gate_173(n244,n94,n242);
and gate_174(n245,n71,n244);
not gate_175(n246,n245);
and gate_176(n247,n237,n246);
and gate_177(n248,n220,n247);
and gate_178(n249,n76,pi6);
not gate_179(n250,n249);
and gate_180(n251,n75,n249);
not gate_181(n252,n251);
and gate_182(n253,n186,n251);
not gate_183(n254,n253);
and gate_184(n255,n248,n254);
not gate_185(po31,n255);
and gate_186(n257,n71,n109);
and gate_187(n258,n71,n184);
not gate_188(n259,n258);
and gate_189(n260,n257,n259);
and gate_190(n261,n134,n260);
not gate_191(n262,n261);
and gate_192(n263,n221,n262);
not gate_193(n264,n263);
and gate_194(n265,n110,n222);
not gate_195(n266,n265);
and gate_196(n267,n213,n266);
not gate_197(n268,n267);
and gate_198(n269,n71,n268);
not gate_199(n270,n269);
and gate_200(n271,n165,n206);
not gate_201(n272,n271);
and gate_202(n273,n270,n272);
not gate_203(n274,n273);
and gate_204(n275,n72,n274);
not gate_205(n276,n275);
and gate_206(n277,n237,n276);
and gate_207(n278,n264,n277);
and gate_208(n279,n71,pi3);
not gate_209(n280,n279);
and gate_210(n281,n203,n280);
not gate_211(n282,n281);
and gate_212(n283,pi3,pi6);
not gate_213(n284,n283);
and gate_214(n285,n74,n77);
not gate_215(n286,n285);
and gate_216(n287,n284,n286);
not gate_217(n288,n287);
and gate_218(n289,n281,n288);
and gate_219(n290,n94,n289);
and gate_220(n291,n184,n290);
not gate_221(n292,n291);
and gate_222(n293,n278,n292);
and gate_223(n294,n190,n196);
not gate_224(n295,n294);
and gate_225(n296,n293,n295);
not gate_226(po32,n296);
and gate_227(n298,n138,n226);
not gate_228(n299,n298);
and gate_229(n300,n75,n77);
not gate_230(n301,n300);
and gate_231(n302,n75,n301);
not gate_232(n303,n302);
and gate_233(n304,pi0,pi2);
not gate_234(n305,n304);
and gate_235(n306,n93,n304);
and gate_236(n307,n302,n306);
and gate_237(n308,n299,n307);
and gate_238(n309,n142,n238);
not gate_239(n310,n309);
and gate_240(n311,n190,n309);
not gate_241(n312,n311);
and gate_242(n313,n308,n312);
not gate_243(po33,n313);
and gate_244(n315,n129,n249);
not gate_245(n316,n315);
and gate_246(n317,n86,n316);
not gate_247(n318,n317);
and gate_248(n319,pi7,n318);
not gate_249(n320,n319);
and gate_250(n321,n146,n199);
not gate_251(n322,n321);
and gate_252(n323,n320,n322);
not gate_253(n324,n323);
and gate_254(n325,n75,n324);
not gate_255(n326,n325);
and gate_256(n327,n129,n167);
not gate_257(n328,n327);
and gate_258(n329,pi1,n76);
not gate_259(n330,n329);
and gate_260(n331,n328,n330);
and gate_261(n332,n86,n250);
not gate_262(n333,n332);
and gate_263(n334,n75,n332);
not gate_264(n335,n334);
and gate_265(n336,n223,n335);
and gate_266(n337,n331,n336);
and gate_267(n338,n326,n337);
and gate_268(n339,n71,n73);
and gate_269(n340,n87,n339);
not gate_270(n341,n340);
and gate_271(n342,n88,n304);
not gate_272(n343,n342);
and gate_273(n344,n341,n343);
not gate_274(n345,n344);
and gate_275(n346,pi6,n345);
not gate_276(n347,n346);
and gate_277(n348,pi2,n77);
and gate_278(n349,pi0,pi4);
and gate_279(n350,n348,n349);
not gate_280(n351,n350);
and gate_281(n352,n347,n351);
not gate_282(n353,n352);
and gate_283(n354,n76,n353);
and gate_284(n355,n72,n354);
not gate_285(n356,n355);
and gate_286(n357,n338,n356);
and gate_287(n358,n74,n85);
not gate_288(n359,n358);
and gate_289(n360,pi3,n249);
and gate_290(n361,n106,n360);
not gate_291(n362,n361);
and gate_292(n363,n359,n362);
not gate_293(n364,n363);
and gate_294(n365,n87,n364);
not gate_295(n366,n365);
and gate_296(n367,n357,n366);
not gate_297(po34,n367);
and gate_298(n369,n72,pi4);
and gate_299(n370,n305,n369);
and gate_300(n371,n71,pi2);
not gate_301(n372,n371);
and gate_302(n373,n166,n372);
not gate_303(n374,n373);
and gate_304(n375,n169,n374);
not gate_305(n376,n375);
and gate_306(n377,n370,n376);
and gate_307(n378,n71,n369);
and gate_308(n379,n74,n76);
not gate_309(n380,n379);
and gate_310(n381,n240,n380);
and gate_311(n382,n378,n381);
not gate_312(n383,n382);
and gate_313(n384,n377,n383);
not gate_314(po35,n384);
and gate_315(n386,n133,n190);
not gate_316(n387,n386);
and gate_317(n388,n71,pi4);
not gate_318(n389,n388);
and gate_319(n390,pi0,n75);
not gate_320(n391,n390);
and gate_321(n392,n389,n391);
not gate_322(n393,n392);
and gate_323(n394,n374,n392);
and gate_324(n395,n72,n76);
not gate_325(n396,n395);
and gate_326(n397,n394,n395);
and gate_327(n398,pi3,n94);
not gate_328(n399,n398);
and gate_329(n400,n183,n399);
not gate_330(n401,n400);
and gate_331(n402,n106,n401);
not gate_332(n403,n402);
and gate_333(n404,n397,n403);
and gate_334(n405,n387,n404);
not gate_335(po36,n405);
and gate_336(n407,pi0,n147);
not gate_337(n408,n407);
and gate_338(n409,n74,n408);
not gate_339(n410,n409);
and gate_340(n411,pi0,n143);
not gate_341(n412,n411);
and gate_342(n413,n175,n412);
not gate_343(n414,n413);
and gate_344(n415,n410,n414);
and gate_345(n416,n72,pi5);
not gate_346(n417,n416);
and gate_347(n418,n330,n417);
not gate_348(n419,n418);
and gate_349(n420,pi0,n419);
not gate_350(n421,n420);
and gate_351(n422,n224,n389);
and gate_352(n423,n421,n422);
and gate_353(n424,pi3,n423);
not gate_354(n425,n424);
and gate_355(n426,n415,n425);
and gate_356(n427,pi1,pi3);
not gate_357(n428,n427);
and gate_358(n429,n72,n74);
not gate_359(n430,n429);
and gate_360(n431,n428,n430);
not gate_361(n432,n431);
and gate_362(n433,n396,n431);
and gate_363(n434,n304,n433);
not gate_364(n435,n434);
and gate_365(n436,n426,n435);
and gate_366(n437,n103,n436);
and gate_367(n438,pi3,n190);
not gate_368(n439,n438);
and gate_369(n440,n437,n439);
not gate_370(po37,n440);
and gate_371(n442,pi0,pi3);
not gate_372(n443,n442);
and gate_373(n444,n71,n74);
not gate_374(n445,n444);
and gate_375(n446,n443,n445);
not gate_376(n447,n446);
and gate_377(n448,n73,n98);
not gate_378(n449,n448);
and gate_379(n450,n447,n448);
and gate_380(n451,n72,n450);
not gate_381(n452,n451);
and gate_382(n453,n239,n392);
not gate_383(n454,n453);
and gate_384(n455,n71,n75);
not gate_385(n456,n455);
and gate_386(n457,n111,n456);
not gate_387(n458,n457);
and gate_388(n459,n454,n458);
not gate_389(n460,n459);
and gate_390(n461,n234,n460);
and gate_391(n462,n452,n461);
and gate_392(n463,n292,n462);
and gate_393(n464,n295,n463);
not gate_394(po38,n464);
and gate_395(n466,n71,n249);
not gate_396(n467,n466);
and gate_397(n468,n75,n467);
and gate_398(n469,n333,n468);
and gate_399(n470,n359,n469);
and gate_400(n471,pi5,n216);
not gate_401(n472,n471);
and gate_402(n473,pi0,n199);
not gate_403(n474,n473);
and gate_404(n475,n472,n474);
not gate_405(n476,n475);
and gate_406(n477,n75,n476);
not gate_407(n478,n477);
and gate_408(n479,n74,n474);
not gate_409(n480,n479);
and gate_410(n481,n477,n480);
not gate_411(n482,n481);
and gate_412(n483,n470,n482);
and gate_413(n484,n142,n190);
not gate_414(n485,n484);
and gate_415(n486,n483,n485);
and gate_416(n487,n146,n204);
not gate_417(n488,n487);
and gate_418(n489,n486,n488);
not gate_419(po39,n489);
and gate_420(n491,n241,n257);
not gate_421(n492,n491);
and gate_422(n493,n221,n492);
not gate_423(n494,n493);
and gate_424(n495,n71,n231);
not gate_425(n496,n495);
and gate_426(n497,pi0,n238);
not gate_427(n498,n497);
and gate_428(n499,n496,n498);
and gate_429(n500,pi2,n280);
not gate_430(n501,n500);
and gate_431(n502,n73,n279);
not gate_432(n503,n502);
and gate_433(n504,n501,n503);
and gate_434(n505,pi1,n504);
not gate_435(n506,n505);
and gate_436(n507,n499,n506);
not gate_437(n508,n507);
and gate_438(n509,n225,n508);
not gate_439(n510,n509);
and gate_440(n511,pi0,n178);
not gate_441(n512,n511);
and gate_442(n513,n129,n210);
not gate_443(n514,n513);
and gate_444(n515,n512,n514);
not gate_445(n516,n515);
and gate_446(n517,pi5,n516);
not gate_447(n518,n517);
and gate_448(n519,n129,n398);
not gate_449(n520,n519);
and gate_450(n521,n518,n520);
not gate_451(n522,n521);
and gate_452(n523,pi2,n522);
not gate_453(n524,n523);
and gate_454(n525,n74,n98);
not gate_455(n526,n525);
and gate_456(n527,n258,n525);
not gate_457(n528,n527);
and gate_458(n529,n524,n528);
and gate_459(n530,n510,n529);
and gate_460(n531,n494,n530);
and gate_461(n532,pi1,n73);
not gate_462(n533,n532);
and gate_463(n534,pi2,pi6);
not gate_464(n535,n534);
and gate_465(n536,n73,n77);
not gate_466(n537,n536);
and gate_467(n538,n535,n537);
not gate_468(n539,n538);
and gate_469(n540,n533,n538);
and gate_470(n541,n239,n540);
and gate_471(n542,pi0,n541);
not gate_472(n543,n542);
and gate_473(n544,n77,n196);
not gate_474(n545,n544);
and gate_475(n546,n543,n545);
not gate_476(n547,n546);
and gate_477(n548,n94,n547);
not gate_478(n549,n548);
and gate_479(n550,n531,n549);
and gate_480(n551,pi2,n78);
and gate_481(n552,pi0,n551);
not gate_482(n553,n552);
and gate_483(n554,pi7,n258);
not gate_484(n555,n554);
and gate_485(n556,n553,n555);
not gate_486(n557,n556);
and gate_487(n558,n123,n249);
not gate_488(n559,n558);
and gate_489(n560,n557,n558);
not gate_490(n561,n560);
and gate_491(n562,n550,n561);
not gate_492(po40,n562);
and gate_493(n564,pi1,n74);
not gate_494(n565,n564);
and gate_495(n566,n72,pi3);
not gate_496(n567,n566);
and gate_497(n568,n565,n567);
not gate_498(n569,n568);
and gate_499(n570,n165,n569);
and gate_500(n571,pi3,n76);
and gate_501(n572,n73,n571);
not gate_502(n573,n572);
and gate_503(n574,n146,n572);
not gate_504(n575,n574);
and gate_505(n576,n570,n575);
not gate_506(po41,n576);
and gate_507(n578,n469,n478);
and gate_508(n579,pi1,n75);
and gate_509(n580,pi0,n579);
and gate_510(n581,n128,n580);
not gate_511(n582,n581);
and gate_512(n583,n578,n582);
and gate_513(n584,n148,n190);
not gate_514(n585,n584);
and gate_515(n586,n583,n585);
not gate_516(po42,n586);
and gate_517(n588,n80,n122);
not gate_518(n589,n588);
and gate_519(n590,n228,n456);
not gate_520(n591,n590);
and gate_521(n592,n589,n591);
not gate_522(n593,n592);
and gate_523(n594,n229,n333);
and gate_524(n595,pi4,n594);
not gate_525(n596,n595);
and gate_526(n597,n71,n329);
not gate_527(n598,n597);
and gate_528(n599,n421,n598);
not gate_529(n600,n599);
and gate_530(n601,n73,n600);
not gate_531(n602,n601);
and gate_532(n603,n174,n602);
not gate_533(n604,n603);
and gate_534(n605,n75,pi6);
and gate_535(n606,n604,n605);
not gate_536(n607,n606);
and gate_537(n608,n596,n607);
and gate_538(n609,n593,n608);
and gate_539(n610,n322,n472);
and gate_540(n611,n142,n551);
not gate_541(n612,n611);
and gate_542(n613,n555,n612);
not gate_543(n614,n613);
and gate_544(n615,n249,n614);
not gate_545(n616,n615);
and gate_546(n617,n610,n616);
not gate_547(n618,n617);
and gate_548(n619,n75,n618);
not gate_549(n620,n619);
and gate_550(n621,n609,n620);
and gate_551(n622,n75,pi7);
not gate_552(n623,n622);
and gate_553(n624,n258,n623);
not gate_554(n625,n624);
and gate_555(n626,n119,n622);
not gate_556(n627,n626);
and gate_557(n628,n625,n627);
not gate_558(n629,n628);
and gate_559(n630,pi6,n629);
not gate_560(n631,n630);
and gate_561(n632,n72,n536);
and gate_562(n633,n388,n632);
not gate_563(n634,n633);
and gate_564(n635,n631,n634);
not gate_565(n636,n635);
and gate_566(n637,n76,n636);
not gate_567(n638,n637);
and gate_568(n639,n73,pi4);
and gate_569(n640,n129,n639);
not gate_570(n641,n640);
and gate_571(n642,pi5,n640);
not gate_572(n643,n642);
and gate_573(n644,n638,n643);
not gate_574(n645,n644);
and gate_575(n646,pi3,n645);
not gate_576(n647,n646);
and gate_577(n648,n106,n178);
not gate_578(n649,n648);
and gate_579(n650,n647,n649);
and gate_580(n651,n621,n650);
not gate_581(po43,n651);
and gate_582(n653,n72,n110);
and gate_583(n654,n393,n653);
and gate_584(n655,n526,n559);
not gate_585(n656,n655);
and gate_586(n657,n186,n656);
not gate_587(n658,n657);
and gate_588(n659,n654,n658);
not gate_589(po44,n659);
and gate_590(n661,n118,n185);
not gate_591(n662,n661);
and gate_592(n663,n71,n641);
and gate_593(n664,n662,n663);
and gate_594(n665,pi5,n662);
not gate_595(n666,n665);
and gate_596(n667,n105,n533);
and gate_597(n668,n76,n667);
and gate_598(n669,n539,n668);
not gate_599(n670,n669);
and gate_600(n671,n666,n670);
not gate_601(n672,n671);
and gate_602(n673,n455,n672);
not gate_603(n674,n673);
and gate_604(n675,n664,n674);
and gate_605(n676,n73,n75);
and gate_606(n677,n199,n676);
and gate_607(n678,n129,n677);
not gate_608(n679,n678);
and gate_609(n680,n675,n679);
not gate_610(po45,n680);
and gate_611(n682,n71,n532);
and gate_612(n683,n525,n682);
not gate_613(n684,n683);
and gate_614(n685,n112,n684);
and gate_615(n686,n201,n685);
not gate_616(po46,n686);
and gate_617(n688,n187,n667);
and gate_618(n689,n120,n259);
not gate_619(n690,n689);
and gate_620(n691,pi4,n690);
not gate_621(n692,n691);
and gate_622(n693,n688,n692);
and gate_623(n694,n71,n665);
not gate_624(n695,n694);
and gate_625(n696,n142,n171);
not gate_626(n697,n696);
and gate_627(n698,n695,n697);
not gate_628(n699,n698);
and gate_629(n700,n75,n699);
not gate_630(n701,n700);
and gate_631(n702,n693,n701);
and gate_632(n703,n71,n669);
not gate_633(n704,n703);
and gate_634(n705,pi2,n85);
not gate_635(n706,n705);
and gate_636(n707,n142,n705);
not gate_637(n708,n707);
and gate_638(n709,n704,n708);
not gate_639(n710,n709);
and gate_640(n711,n75,n710);
not gate_641(n712,n711);
and gate_642(n713,n702,n712);
and gate_643(n714,n126,n713);
and gate_644(n715,pi2,n193);
and gate_645(n716,n142,n715);
not gate_646(n717,n716);
and gate_647(n718,n73,n76);
not gate_648(n719,n718);
and gate_649(n720,n129,n718);
not gate_650(n721,n720);
and gate_651(n722,n717,n721);
not gate_652(n723,n722);
and gate_653(n724,n92,n723);
and gate_654(n725,n75,n724);
not gate_655(n726,n725);
and gate_656(n727,n714,n726);
not gate_657(po47,n727);
and gate_658(n729,n75,n588);
not gate_659(n730,n729);
and gate_660(n731,n129,n151);
and gate_661(n732,n101,n731);
and gate_662(n733,n730,n732);
not gate_663(po48,n733);
and gate_664(n735,pi2,pi4);
and gate_665(n736,n129,n735);
not gate_666(n737,n736);
and gate_667(n738,pi3,n736);
not gate_668(n739,n738);
and gate_669(n740,n260,n739);
and gate_670(n741,n99,n252);
not gate_671(n742,n741);
and gate_672(n743,n106,n742);
not gate_673(n744,n743);
and gate_674(n745,n740,n744);
not gate_675(po49,n745);
and gate_676(n747,n128,n676);
and gate_677(n748,n192,n747);
and gate_678(n749,n144,n190);
not gate_679(n750,n749);
and gate_680(n751,n748,n750);
not gate_681(po50,n751);
and gate_682(n753,n109,n147);
and gate_683(n754,n737,n753);
and gate_684(n755,n120,n130);
not gate_685(n756,n755);
and gate_686(n757,n98,n756);
not gate_687(n758,n757);
and gate_688(n759,n754,n758);
and gate_689(n760,pi0,n427);
not gate_690(n761,n760);
and gate_691(n762,n179,n207);
not gate_692(n763,n762);
and gate_693(n764,n129,n763);
not gate_694(n765,n764);
and gate_695(n766,n761,n765);
not gate_696(n767,n766);
and gate_697(n768,n73,n767);
not gate_698(n769,n768);
and gate_699(n770,n106,n206);
not gate_700(n771,n770);
and gate_701(n772,n769,n771);
and gate_702(n773,n759,n772);
and gate_703(n774,pi0,n532);
and gate_704(n775,n358,n774);
not gate_705(n776,n775);
and gate_706(n777,n71,n566);
not gate_707(n778,n777);
and gate_708(n779,pi0,n564);
not gate_709(n780,n779);
and gate_710(n781,n778,n780);
and gate_711(n782,n310,n781);
not gate_712(n783,n782);
and gate_713(n784,n249,n783);
not gate_714(n785,n784);
and gate_715(n786,n776,n785);
not gate_716(n787,n786);
and gate_717(n788,n75,n787);
not gate_718(n789,n788);
and gate_719(n790,n773,n789);
and gate_720(n791,po05,n144);
not gate_721(n792,n791);
and gate_722(n793,n790,n792);
not gate_723(po51,n793);
and gate_724(n795,n73,n206);
not gate_725(n796,n795);
and gate_726(n797,pi4,n230);
and gate_727(n798,n443,n797);
not gate_728(n799,n798);
and gate_729(n800,n796,n799);
not gate_730(n801,n800);
and gate_731(n802,n72,n801);
not gate_732(n803,n802);
and gate_733(n804,n109,n443);
and gate_734(n805,n99,n804);
and gate_735(n806,n803,n805);
and gate_736(n807,n72,n131);
not gate_737(n808,n807);
and gate_738(n809,n781,n808);
not gate_739(n810,n809);
and gate_740(n811,n251,n810);
not gate_741(n812,n811);
and gate_742(n813,n806,n812);
not gate_743(po52,n813);
and gate_744(n815,pi1,n110);
not gate_745(n816,n815);
and gate_746(n817,n243,n816);
not gate_747(n818,n817);
and gate_748(n819,n76,n818);
not gate_749(n820,n819);
and gate_750(n821,pi5,n231);
and gate_751(n822,pi1,n821);
not gate_752(n823,n822);
and gate_753(n824,n820,n823);
not gate_754(n825,n824);
and gate_755(n826,n75,n825);
not gate_756(n827,n826);
and gate_757(n828,n75,n230);
not gate_758(n829,n828);
and gate_759(n830,pi1,n111);
not gate_760(n831,n830);
and gate_761(n832,n829,n831);
not gate_762(n833,n832);
and gate_763(n834,n827,n833);
and gate_764(n835,n282,n526);
and gate_765(n836,pi2,n835);
not gate_766(n837,n836);
and gate_767(n838,n165,n525);
not gate_768(n839,n838);
and gate_769(n840,n837,n839);
not gate_770(n841,n840);
and gate_771(n842,pi1,n841);
not gate_772(n843,n842);
and gate_773(n844,n159,n226);
not gate_774(n845,n844);
and gate_775(n846,n843,n845);
and gate_776(n847,n834,n846);
and gate_777(n848,n231,n249);
and gate_778(n849,pi1,n848);
not gate_779(n850,n849);
and gate_780(n851,n85,n818);
not gate_781(n852,n851);
and gate_782(n853,n850,n852);
not gate_783(n854,n853);
and gate_784(n855,n71,n854);
not gate_785(n856,n855);
and gate_786(n857,n184,n358);
not gate_787(n858,n857);
and gate_788(n859,n250,n706);
not gate_789(n860,n859);
and gate_790(n861,n427,n860);
not gate_791(n862,n861);
and gate_792(n863,n858,n862);
not gate_793(n864,n863);
and gate_794(n865,pi0,n864);
not gate_795(n866,n865);
and gate_796(n867,n856,n866);
not gate_797(n868,n867);
and gate_798(n869,n75,n868);
not gate_799(n870,n869);
and gate_800(n871,n847,n870);
and gate_801(n872,n71,n818);
not gate_802(n873,n872);
and gate_803(n874,pi0,n568);
and gate_804(n875,n241,n874);
not gate_805(n876,n875);
and gate_806(n877,n873,n876);
not gate_807(n878,n877);
and gate_808(n879,po05,n878);
not gate_809(n880,n879);
and gate_810(n881,n871,n880);
not gate_811(po53,n881);
and gate_812(n883,n243,n310);
and gate_813(n884,n179,n211);
not gate_814(n885,n884);
and gate_815(n886,n774,n885);
not gate_816(n887,n886);
and gate_817(n888,n883,n887);
and gate_818(n889,n75,n147);
not gate_819(n890,n889);
and gate_820(n891,n231,n890);
not gate_821(n892,n891);
and gate_822(n893,n888,n892);
and gate_823(n894,n74,pi5);
and gate_824(n895,n73,n894);
not gate_825(n896,n895);
and gate_826(n897,n108,n895);
not gate_827(n898,n897);
and gate_828(n899,n496,n780);
not gate_829(n900,n899);
and gate_830(n901,n76,n900);
not gate_831(n902,n901);
and gate_832(n903,n898,n902);
not gate_833(n904,n903);
and gate_834(n905,n75,n904);
not gate_835(n906,n905);
and gate_836(n907,n893,n906);
and gate_837(n908,n71,n131);
not gate_838(n909,n908);
and gate_839(n910,n281,n909);
not gate_840(n911,n910);
and gate_841(n912,n85,n911);
not gate_842(n913,n912);
and gate_843(n914,n241,n466);
not gate_844(n915,n914);
and gate_845(n916,n913,n915);
not gate_846(n917,n916);
and gate_847(n918,pi1,n917);
not gate_848(n919,n918);
and gate_849(n920,n85,n232);
not gate_850(n921,n920);
and gate_851(n922,n919,n921);
not gate_852(n923,n922);
and gate_853(n924,n75,n923);
not gate_854(n925,n924);
and gate_855(n926,n907,n925);
and gate_856(n927,pi1,n911);
not gate_857(n928,n927);
and gate_858(n929,n233,n928);
not gate_859(n930,n929);
and gate_860(n931,po05,n930);
not gate_861(n932,n931);
and gate_862(n933,n926,n932);
not gate_863(po54,n933);
and gate_864(n935,n98,n108);
not gate_865(n936,n935);
and gate_866(n937,pi1,n936);
and gate_867(n938,n75,n95);
not gate_868(n939,n938);
and gate_869(n940,pi2,n939);
not gate_870(n941,n940);
and gate_871(n942,n449,n941);
not gate_872(n943,n942);
and gate_873(n944,n142,n943);
not gate_874(n945,n944);
and gate_875(n946,n937,n945);
and gate_876(n947,n249,n305);
not gate_877(n948,n947);
and gate_878(n949,pi0,n705);
not gate_879(n950,n949);
and gate_880(n951,n948,n950);
not gate_881(n952,n951);
and gate_882(n953,n579,n952);
not gate_883(n954,n953);
and gate_884(n955,n946,n954);
and gate_885(n956,n75,n82);
not gate_886(n957,n956);
and gate_887(n958,n144,n957);
not gate_888(n959,n958);
and gate_889(n960,n955,n959);
and gate_890(n961,po05,n119);
not gate_891(n962,n961);
and gate_892(n963,n960,n962);
not gate_893(po55,n963);
and gate_894(n965,n71,n735);
not gate_895(n966,n965);
and gate_896(n967,n104,n210);
not gate_897(n968,n967);
and gate_898(n969,n816,n968);
and gate_899(n970,n966,n969);
and gate_900(n971,n71,n259);
and gate_901(n972,n970,n971);
and gate_902(n973,pi2,pi5);
not gate_903(n974,n973);
and gate_904(n975,n719,n974);
and gate_905(n976,n111,n975);
and gate_906(n977,n567,n976);
and gate_907(n978,n455,n977);
not gate_908(n979,n978);
and gate_909(n980,n972,n979);
and gate_910(n981,n567,n705);
and gate_911(n982,n455,n981);
not gate_912(n983,n982);
and gate_913(n984,n980,n983);
and gate_914(n985,n573,n974);
not gate_915(n986,n985);
and gate_916(n987,n567,n986);
and gate_917(n988,n92,n987);
and gate_918(n989,n455,n988);
not gate_919(n990,n989);
and gate_920(n991,n984,n990);
not gate_921(po56,n991);
and gate_922(n993,n282,n532);
not gate_923(n994,n993);
and gate_924(n995,n136,n994);
and gate_925(n996,n147,n966);
and gate_926(n997,n689,n996);
and gate_927(n998,n995,n997);
and gate_928(n999,n172,n896);
not gate_929(n1000,n999);
and gate_930(n1001,n71,n1000);
not gate_931(n1002,n1001);
and gate_932(n1003,n165,n193);
not gate_933(n1004,n1003);
and gate_934(n1005,n1002,n1004);
not gate_935(n1006,n1005);
and gate_936(n1007,pi1,n1006);
not gate_937(n1008,n1007);
and gate_938(n1009,n106,n571);
not gate_939(n1010,n1009);
and gate_940(n1011,n1008,n1010);
not gate_941(n1012,n1011);
and gate_942(n1013,n75,n1012);
not gate_943(n1014,n1013);
and gate_944(n1015,n998,n1014);
and gate_945(n1016,n430,n705);
and gate_946(n1017,n455,n1016);
not gate_947(n1018,n1017);
and gate_948(n1019,n1015,n1018);
and gate_949(n1020,n73,n379);
not gate_950(n1021,n1020);
and gate_951(n1022,n974,n1021);
not gate_952(n1023,n1022);
and gate_953(n1024,n71,n1023);
not gate_954(n1025,n1024);
and gate_955(n1026,n165,n571);
not gate_956(n1027,n1026);
and gate_957(n1028,n1025,n1027);
not gate_958(n1029,n1028);
and gate_959(n1030,pi1,n1029);
not gate_960(n1031,n1030);
and gate_961(n1032,n129,n715);
not gate_962(n1033,n1032);
and gate_963(n1034,n1031,n1033);
not gate_964(n1035,n1034);
and gate_965(n1036,n92,n1035);
and gate_966(n1037,n75,n1036);
not gate_967(n1038,n1037);
and gate_968(n1039,n1019,n1038);
not gate_969(po57,n1039);
and gate_970(n1041,pi3,n156);
and gate_971(n1042,n662,n692);
and gate_972(n1043,n701,n1042);
and gate_973(n1044,n712,n1043);
and gate_974(n1045,n1041,n1044);
and gate_975(n1046,n142,n973);
not gate_976(n1047,n1046);
and gate_977(n1048,n721,n1047);
not gate_978(n1049,n1048);
and gate_979(n1050,n92,n1049);
and gate_980(n1051,n210,n1050);
not gate_981(n1052,n1051);
and gate_982(n1053,n1045,n1052);
not gate_983(po58,n1053);
and gate_984(n1055,pi4,n305);
not gate_985(n1056,n1055);
and gate_986(n1057,n99,n1056);
and gate_987(n1058,pi0,n539);
not gate_988(n1059,n1058);
and gate_989(n1060,n71,n77);
not gate_990(n1061,n1060);
and gate_991(n1062,n1059,n1061);
not gate_992(n1063,n1062);
and gate_993(n1064,n94,n1063);
not gate_994(n1065,n1064);
and gate_995(n1066,n1057,n1065);
and gate_996(n1067,n140,n187);
not gate_997(n1068,n1067);
and gate_998(n1069,n251,n1068);
not gate_999(n1070,n1069);
and gate_1000(n1071,n1066,n1070);
and gate_1001(n1072,n303,n432);
and gate_1002(n1073,pi2,n1072);
not gate_1003(n1074,n1073);
and gate_1004(n1075,n605,n815);
not gate_1005(n1076,n1075);
and gate_1006(n1077,n1074,n1076);
not gate_1007(n1078,n1077);
and gate_1008(n1079,n76,n1078);
not gate_1009(n1080,n1079);
and gate_1010(n1081,n222,n432);
and gate_1011(n1082,pi2,n1081);
not gate_1012(n1083,n1082);
and gate_1013(n1084,n1080,n1083);
not gate_1014(n1085,n1084);
and gate_1015(n1086,pi0,n1085);
not gate_1016(n1087,n1086);
and gate_1017(n1088,n210,n249);
not gate_1018(n1089,n1088);
and gate_1019(n1090,n106,n1088);
not gate_1020(n1091,n1090);
and gate_1021(n1092,n1087,n1091);
and gate_1022(n1093,n1071,n1092);
and gate_1023(n1094,pi2,n808);
not gate_1024(n1095,n1094);
and gate_1025(n1096,n71,n1095);
not gate_1026(n1097,n1096);
and gate_1027(n1098,n163,n1097);
not gate_1028(n1099,n1098);
and gate_1029(n1100,n96,n1099);
not gate_1030(n1101,n1100);
and gate_1031(n1102,n1093,n1101);
not gate_1032(po59,n1102);
and gate_1033(n1104,n392,n753);
and gate_1034(n1105,n443,n1104);
and gate_1035(n1106,n75,n232);
not gate_1036(n1107,n1106);
and gate_1037(n1108,n1105,n1107);
and gate_1038(n1109,n246,n1108);
and gate_1039(n1110,n85,n242);
and gate_1040(n1111,n455,n1110);
not gate_1041(n1112,n1111);
and gate_1042(n1113,n1109,n1112);
and gate_1043(n1114,po05,n242);
and gate_1044(n1115,n71,n1114);
not gate_1045(n1116,n1115);
and gate_1046(n1117,n1113,n1116);
not gate_1047(po60,n1117);
and gate_1048(n1119,n226,n1089);
and gate_1049(n1120,n149,n845);
and gate_1050(n1121,n1119,n1120);
not gate_1051(po61,n1121);
and gate_1052(n1123,n252,n779);
and gate_1053(n1124,n526,n1123);
not gate_1054(po62,n1124);
endmodule
